* SPICE3 file created from attempt3.ext - technology: scmos

.option scale=0.3u

M1000 attempt2_4/OR2X1_1/a_9_54# attempt2_4/m1_133_n102# attempt2_4/OR2X1_1/a_2_54# attempt2_4/OR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1001 attempt2_4/OR2X1_1/vdd attempt2_4/Input2 attempt2_4/OR2X1_1/a_9_54# attempt2_4/OR2X1_1/vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1002 attempt2_4/Output2 attempt2_4/OR2X1_1/a_2_54# attempt2_4/OR2X1_1/vdd attempt2_4/OR2X1_1/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1003 attempt2_4/OR2X1_1/a_2_54# attempt2_4/m1_133_n102# attempt2_4/OR2X1_1/gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=110 ps=62
M1004 attempt2_4/OR2X1_1/gnd attempt2_4/Input2 attempt2_4/OR2X1_1/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 attempt2_4/Output2 attempt2_4/OR2X1_1/a_2_54# attempt2_4/OR2X1_1/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1006 attempt2_4/XOR2X1_1/vdd attempt2_4/m1_n54_n42# attempt2_4/XOR2X1_1/a_2_6# attempt2_4/XOR2X1_1/vdd pfet w=40 l=2
+  ad=560 pd=188 as=200 ps=90
M1007 attempt2_4/XOR2X1_1/a_18_54# attempt2_4/XOR2X1_1/a_13_43# attempt2_4/XOR2X1_1/vdd attempt2_4/XOR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1008 attempt2_4/m1_133_n102# attempt2_4/m1_n54_n42# attempt2_4/XOR2X1_1/a_18_54# attempt2_4/XOR2X1_1/vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1009 attempt2_4/XOR2X1_1/a_35_54# attempt2_4/XOR2X1_1/a_2_6# attempt2_4/m1_133_n102# attempt2_4/XOR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1010 attempt2_4/XOR2X1_1/vdd attempt2_4/m1_71_n159# attempt2_4/XOR2X1_1/a_35_54# attempt2_4/XOR2X1_1/vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 attempt2_4/XOR2X1_1/a_13_43# attempt2_4/m1_71_n159# attempt2_4/XOR2X1_1/vdd attempt2_4/XOR2X1_1/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1012 attempt2_4/XOR2X1_1/gnd attempt2_4/m1_n54_n42# attempt2_4/XOR2X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=280 pd=108 as=100 ps=50
M1013 attempt2_4/XOR2X1_1/a_18_6# attempt2_4/XOR2X1_1/a_13_43# attempt2_4/XOR2X1_1/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1014 attempt2_4/m1_133_n102# attempt2_4/XOR2X1_1/a_2_6# attempt2_4/XOR2X1_1/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1015 attempt2_4/XOR2X1_1/a_35_6# attempt2_4/m1_n54_n42# attempt2_4/m1_133_n102# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1016 attempt2_4/XOR2X1_1/gnd attempt2_4/m1_71_n159# attempt2_4/XOR2X1_1/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1017 attempt2_4/XOR2X1_1/a_13_43# attempt2_4/m1_71_n159# attempt2_4/XOR2X1_1/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1018 attempt2_4/DFFPOSX1_2/vdd attempt2_4/m1_n35_n168# attempt2_4/DFFPOSX1_2/a_2_6# attempt2_4/DFFPOSX1_2/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1019 attempt2_4/DFFPOSX1_2/a_17_74# attempt2_4/m1_n64_n214# attempt2_4/DFFPOSX1_2/vdd attempt2_4/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1020 attempt2_4/DFFPOSX1_2/a_22_6# attempt2_4/m1_n35_n168# attempt2_4/DFFPOSX1_2/a_17_74# attempt2_4/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1021 attempt2_4/DFFPOSX1_2/a_31_74# attempt2_4/DFFPOSX1_2/a_2_6# attempt2_4/DFFPOSX1_2/a_22_6# attempt2_4/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1022 attempt2_4/DFFPOSX1_2/vdd attempt2_4/DFFPOSX1_2/a_34_4# attempt2_4/DFFPOSX1_2/a_31_74# attempt2_4/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1023 attempt2_4/DFFPOSX1_2/a_34_4# attempt2_4/DFFPOSX1_2/a_22_6# attempt2_4/DFFPOSX1_2/vdd attempt2_4/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1024 attempt2_4/DFFPOSX1_2/a_61_74# attempt2_4/DFFPOSX1_2/a_34_4# attempt2_4/DFFPOSX1_2/vdd attempt2_4/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1025 attempt2_4/DFFPOSX1_2/a_66_6# attempt2_4/DFFPOSX1_2/a_2_6# attempt2_4/DFFPOSX1_2/a_61_74# attempt2_4/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1026 attempt2_4/DFFPOSX1_2/a_76_84# attempt2_4/m1_n35_n168# attempt2_4/DFFPOSX1_2/a_66_6# attempt2_4/DFFPOSX1_2/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1027 attempt2_4/DFFPOSX1_2/vdd attempt2_4/m1_71_n159# attempt2_4/DFFPOSX1_2/a_76_84# attempt2_4/DFFPOSX1_2/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 attempt2_4/DFFPOSX1_2/gnd attempt2_4/m1_n35_n168# attempt2_4/DFFPOSX1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1029 attempt2_4/m1_71_n159# attempt2_4/DFFPOSX1_2/a_66_6# attempt2_4/DFFPOSX1_2/vdd attempt2_4/DFFPOSX1_2/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1030 attempt2_4/DFFPOSX1_2/a_17_6# attempt2_4/m1_n64_n214# attempt2_4/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1031 attempt2_4/DFFPOSX1_2/a_22_6# attempt2_4/DFFPOSX1_2/a_2_6# attempt2_4/DFFPOSX1_2/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1032 attempt2_4/DFFPOSX1_2/a_31_6# attempt2_4/m1_n35_n168# attempt2_4/DFFPOSX1_2/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1033 attempt2_4/DFFPOSX1_2/gnd attempt2_4/DFFPOSX1_2/a_34_4# attempt2_4/DFFPOSX1_2/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1034 attempt2_4/DFFPOSX1_2/a_34_4# attempt2_4/DFFPOSX1_2/a_22_6# attempt2_4/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1035 attempt2_4/DFFPOSX1_2/a_61_6# attempt2_4/DFFPOSX1_2/a_34_4# attempt2_4/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1036 attempt2_4/DFFPOSX1_2/a_66_6# attempt2_4/m1_n35_n168# attempt2_4/DFFPOSX1_2/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1037 attempt2_4/DFFPOSX1_2/a_76_6# attempt2_4/DFFPOSX1_2/a_2_6# attempt2_4/DFFPOSX1_2/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1038 attempt2_4/DFFPOSX1_2/gnd attempt2_4/m1_71_n159# attempt2_4/DFFPOSX1_2/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1039 attempt2_4/m1_71_n159# attempt2_4/DFFPOSX1_2/a_66_6# attempt2_4/DFFPOSX1_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1040 attempt2_4/OR2X1_0/a_9_54# attempt2_4/Input3 attempt2_4/OR2X1_0/a_2_54# attempt2_4/OR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1041 attempt2_4/OR2X1_0/vdd attempt2_4/m1_133_15# attempt2_4/OR2X1_0/a_9_54# attempt2_4/OR2X1_0/vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1042 attempt2_4/Output1 attempt2_4/OR2X1_0/a_2_54# attempt2_4/OR2X1_0/vdd attempt2_4/OR2X1_0/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1043 attempt2_4/OR2X1_0/a_2_54# attempt2_4/Input3 attempt2_4/OR2X1_0/gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=110 ps=62
M1044 attempt2_4/OR2X1_0/gnd attempt2_4/m1_133_15# attempt2_4/OR2X1_0/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1045 attempt2_4/Output1 attempt2_4/OR2X1_0/a_2_54# attempt2_4/OR2X1_0/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1046 attempt2_4/XOR2X1_0/vdd attempt2_4/m1_n54_n42# attempt2_4/XOR2X1_0/a_2_6# attempt2_4/XOR2X1_0/vdd pfet w=40 l=2
+  ad=560 pd=188 as=200 ps=90
M1047 attempt2_4/XOR2X1_0/a_18_54# attempt2_4/XOR2X1_0/a_13_43# attempt2_4/XOR2X1_0/vdd attempt2_4/XOR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1048 attempt2_4/m1_133_15# attempt2_4/m1_n54_n42# attempt2_4/XOR2X1_0/a_18_54# attempt2_4/XOR2X1_0/vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1049 attempt2_4/XOR2X1_0/a_35_54# attempt2_4/XOR2X1_0/a_2_6# attempt2_4/m1_133_15# attempt2_4/XOR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1050 attempt2_4/XOR2X1_0/vdd attempt2_4/m1_n64_n214# attempt2_4/XOR2X1_0/a_35_54# attempt2_4/XOR2X1_0/vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1051 attempt2_4/XOR2X1_0/a_13_43# attempt2_4/m1_n64_n214# attempt2_4/XOR2X1_0/vdd attempt2_4/XOR2X1_0/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1052 attempt2_4/XOR2X1_0/gnd attempt2_4/m1_n54_n42# attempt2_4/XOR2X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=280 pd=108 as=100 ps=50
M1053 attempt2_4/XOR2X1_0/a_18_6# attempt2_4/XOR2X1_0/a_13_43# attempt2_4/XOR2X1_0/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1054 attempt2_4/m1_133_15# attempt2_4/XOR2X1_0/a_2_6# attempt2_4/XOR2X1_0/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1055 attempt2_4/XOR2X1_0/a_35_6# attempt2_4/m1_n54_n42# attempt2_4/m1_133_15# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1056 attempt2_4/XOR2X1_0/gnd attempt2_4/m1_n64_n214# attempt2_4/XOR2X1_0/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1057 attempt2_4/XOR2X1_0/a_13_43# attempt2_4/m1_n64_n214# attempt2_4/XOR2X1_0/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1058 attempt2_4/DFFPOSX1_1/vdd attempt2_4/m1_n31_n51# attempt2_4/DFFPOSX1_1/a_2_6# attempt2_4/DFFPOSX1_1/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1059 attempt2_4/DFFPOSX1_1/a_17_74# attempt2_4/m1_n54_n42# attempt2_4/DFFPOSX1_1/vdd attempt2_4/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1060 attempt2_4/DFFPOSX1_1/a_22_6# attempt2_4/m1_n31_n51# attempt2_4/DFFPOSX1_1/a_17_74# attempt2_4/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1061 attempt2_4/DFFPOSX1_1/a_31_74# attempt2_4/DFFPOSX1_1/a_2_6# attempt2_4/DFFPOSX1_1/a_22_6# attempt2_4/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1062 attempt2_4/DFFPOSX1_1/vdd attempt2_4/DFFPOSX1_1/a_34_4# attempt2_4/DFFPOSX1_1/a_31_74# attempt2_4/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 attempt2_4/DFFPOSX1_1/a_34_4# attempt2_4/DFFPOSX1_1/a_22_6# attempt2_4/DFFPOSX1_1/vdd attempt2_4/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1064 attempt2_4/DFFPOSX1_1/a_61_74# attempt2_4/DFFPOSX1_1/a_34_4# attempt2_4/DFFPOSX1_1/vdd attempt2_4/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1065 attempt2_4/DFFPOSX1_1/a_66_6# attempt2_4/DFFPOSX1_1/a_2_6# attempt2_4/DFFPOSX1_1/a_61_74# attempt2_4/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1066 attempt2_4/DFFPOSX1_1/a_76_84# attempt2_4/m1_n31_n51# attempt2_4/DFFPOSX1_1/a_66_6# attempt2_4/DFFPOSX1_1/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1067 attempt2_4/DFFPOSX1_1/vdd attempt2_4/m1_n64_n214# attempt2_4/DFFPOSX1_1/a_76_84# attempt2_4/DFFPOSX1_1/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1068 attempt2_4/DFFPOSX1_1/gnd attempt2_4/m1_n31_n51# attempt2_4/DFFPOSX1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1069 attempt2_4/m1_n64_n214# attempt2_4/DFFPOSX1_1/a_66_6# attempt2_4/DFFPOSX1_1/vdd attempt2_4/DFFPOSX1_1/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1070 attempt2_4/DFFPOSX1_1/a_17_6# attempt2_4/m1_n54_n42# attempt2_4/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1071 attempt2_4/DFFPOSX1_1/a_22_6# attempt2_4/DFFPOSX1_1/a_2_6# attempt2_4/DFFPOSX1_1/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1072 attempt2_4/DFFPOSX1_1/a_31_6# attempt2_4/m1_n31_n51# attempt2_4/DFFPOSX1_1/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1073 attempt2_4/DFFPOSX1_1/gnd attempt2_4/DFFPOSX1_1/a_34_4# attempt2_4/DFFPOSX1_1/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1074 attempt2_4/DFFPOSX1_1/a_34_4# attempt2_4/DFFPOSX1_1/a_22_6# attempt2_4/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1075 attempt2_4/DFFPOSX1_1/a_61_6# attempt2_4/DFFPOSX1_1/a_34_4# attempt2_4/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1076 attempt2_4/DFFPOSX1_1/a_66_6# attempt2_4/m1_n31_n51# attempt2_4/DFFPOSX1_1/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1077 attempt2_4/DFFPOSX1_1/a_76_6# attempt2_4/DFFPOSX1_1/a_2_6# attempt2_4/DFFPOSX1_1/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1078 attempt2_4/DFFPOSX1_1/gnd attempt2_4/m1_n64_n214# attempt2_4/DFFPOSX1_1/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1079 attempt2_4/m1_n64_n214# attempt2_4/DFFPOSX1_1/a_66_6# attempt2_4/DFFPOSX1_1/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1080 attempt2_4/DFFPOSX1_0/vdd attempt2_4/m1_n29_66# attempt2_4/DFFPOSX1_0/a_2_6# attempt2_4/DFFPOSX1_0/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1081 attempt2_4/DFFPOSX1_0/a_17_74# attempt2_4/Input1 attempt2_4/DFFPOSX1_0/vdd attempt2_4/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1082 attempt2_4/DFFPOSX1_0/a_22_6# attempt2_4/m1_n29_66# attempt2_4/DFFPOSX1_0/a_17_74# attempt2_4/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1083 attempt2_4/DFFPOSX1_0/a_31_74# attempt2_4/DFFPOSX1_0/a_2_6# attempt2_4/DFFPOSX1_0/a_22_6# attempt2_4/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1084 attempt2_4/DFFPOSX1_0/vdd attempt2_4/DFFPOSX1_0/a_34_4# attempt2_4/DFFPOSX1_0/a_31_74# attempt2_4/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1085 attempt2_4/DFFPOSX1_0/a_34_4# attempt2_4/DFFPOSX1_0/a_22_6# attempt2_4/DFFPOSX1_0/vdd attempt2_4/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1086 attempt2_4/DFFPOSX1_0/a_61_74# attempt2_4/DFFPOSX1_0/a_34_4# attempt2_4/DFFPOSX1_0/vdd attempt2_4/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1087 attempt2_4/DFFPOSX1_0/a_66_6# attempt2_4/DFFPOSX1_0/a_2_6# attempt2_4/DFFPOSX1_0/a_61_74# attempt2_4/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1088 attempt2_4/DFFPOSX1_0/a_76_84# attempt2_4/m1_n29_66# attempt2_4/DFFPOSX1_0/a_66_6# attempt2_4/DFFPOSX1_0/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1089 attempt2_4/DFFPOSX1_0/vdd attempt2_4/m1_n54_n42# attempt2_4/DFFPOSX1_0/a_76_84# attempt2_4/DFFPOSX1_0/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1090 attempt2_4/DFFPOSX1_0/gnd attempt2_4/m1_n29_66# attempt2_4/DFFPOSX1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1091 attempt2_4/m1_n54_n42# attempt2_4/DFFPOSX1_0/a_66_6# attempt2_4/DFFPOSX1_0/vdd attempt2_4/DFFPOSX1_0/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1092 attempt2_4/DFFPOSX1_0/a_17_6# attempt2_4/Input1 attempt2_4/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1093 attempt2_4/DFFPOSX1_0/a_22_6# attempt2_4/DFFPOSX1_0/a_2_6# attempt2_4/DFFPOSX1_0/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1094 attempt2_4/DFFPOSX1_0/a_31_6# attempt2_4/m1_n29_66# attempt2_4/DFFPOSX1_0/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1095 attempt2_4/DFFPOSX1_0/gnd attempt2_4/DFFPOSX1_0/a_34_4# attempt2_4/DFFPOSX1_0/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1096 attempt2_4/DFFPOSX1_0/a_34_4# attempt2_4/DFFPOSX1_0/a_22_6# attempt2_4/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1097 attempt2_4/DFFPOSX1_0/a_61_6# attempt2_4/DFFPOSX1_0/a_34_4# attempt2_4/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1098 attempt2_4/DFFPOSX1_0/a_66_6# attempt2_4/m1_n29_66# attempt2_4/DFFPOSX1_0/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1099 attempt2_4/DFFPOSX1_0/a_76_6# attempt2_4/DFFPOSX1_0/a_2_6# attempt2_4/DFFPOSX1_0/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1100 attempt2_4/DFFPOSX1_0/gnd attempt2_4/m1_n54_n42# attempt2_4/DFFPOSX1_0/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 attempt2_4/m1_n54_n42# attempt2_4/DFFPOSX1_0/a_66_6# attempt2_4/DFFPOSX1_0/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1102 attempt2_3/OR2X1_1/a_9_54# attempt2_3/m1_133_n102# attempt2_3/OR2X1_1/a_2_54# attempt2_3/OR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1103 attempt2_3/OR2X1_1/vdd attempt2_3/Input2 attempt2_3/OR2X1_1/a_9_54# attempt2_3/OR2X1_1/vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1104 attempt2_4/Input2 attempt2_3/OR2X1_1/a_2_54# attempt2_3/OR2X1_1/vdd attempt2_3/OR2X1_1/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1105 attempt2_3/OR2X1_1/a_2_54# attempt2_3/m1_133_n102# attempt2_3/OR2X1_1/gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=110 ps=62
M1106 attempt2_3/OR2X1_1/gnd attempt2_3/Input2 attempt2_3/OR2X1_1/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1107 attempt2_4/Input2 attempt2_3/OR2X1_1/a_2_54# attempt2_3/OR2X1_1/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1108 attempt2_3/XOR2X1_1/vdd attempt2_3/m1_n54_n42# attempt2_3/XOR2X1_1/a_2_6# attempt2_3/XOR2X1_1/vdd pfet w=40 l=2
+  ad=560 pd=188 as=200 ps=90
M1109 attempt2_3/XOR2X1_1/a_18_54# attempt2_3/XOR2X1_1/a_13_43# attempt2_3/XOR2X1_1/vdd attempt2_3/XOR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1110 attempt2_3/m1_133_n102# attempt2_3/m1_n54_n42# attempt2_3/XOR2X1_1/a_18_54# attempt2_3/XOR2X1_1/vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1111 attempt2_3/XOR2X1_1/a_35_54# attempt2_3/XOR2X1_1/a_2_6# attempt2_3/m1_133_n102# attempt2_3/XOR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1112 attempt2_3/XOR2X1_1/vdd attempt2_3/m1_71_n159# attempt2_3/XOR2X1_1/a_35_54# attempt2_3/XOR2X1_1/vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1113 attempt2_3/XOR2X1_1/a_13_43# attempt2_3/m1_71_n159# attempt2_3/XOR2X1_1/vdd attempt2_3/XOR2X1_1/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1114 attempt2_3/XOR2X1_1/gnd attempt2_3/m1_n54_n42# attempt2_3/XOR2X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=280 pd=108 as=100 ps=50
M1115 attempt2_3/XOR2X1_1/a_18_6# attempt2_3/XOR2X1_1/a_13_43# attempt2_3/XOR2X1_1/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1116 attempt2_3/m1_133_n102# attempt2_3/XOR2X1_1/a_2_6# attempt2_3/XOR2X1_1/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1117 attempt2_3/XOR2X1_1/a_35_6# attempt2_3/m1_n54_n42# attempt2_3/m1_133_n102# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1118 attempt2_3/XOR2X1_1/gnd attempt2_3/m1_71_n159# attempt2_3/XOR2X1_1/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1119 attempt2_3/XOR2X1_1/a_13_43# attempt2_3/m1_71_n159# attempt2_3/XOR2X1_1/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1120 attempt2_3/DFFPOSX1_2/vdd attempt2_3/m1_n35_n168# attempt2_3/DFFPOSX1_2/a_2_6# attempt2_3/DFFPOSX1_2/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1121 attempt2_3/DFFPOSX1_2/a_17_74# attempt2_3/m1_n64_n214# attempt2_3/DFFPOSX1_2/vdd attempt2_3/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1122 attempt2_3/DFFPOSX1_2/a_22_6# attempt2_3/m1_n35_n168# attempt2_3/DFFPOSX1_2/a_17_74# attempt2_3/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1123 attempt2_3/DFFPOSX1_2/a_31_74# attempt2_3/DFFPOSX1_2/a_2_6# attempt2_3/DFFPOSX1_2/a_22_6# attempt2_3/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1124 attempt2_3/DFFPOSX1_2/vdd attempt2_3/DFFPOSX1_2/a_34_4# attempt2_3/DFFPOSX1_2/a_31_74# attempt2_3/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1125 attempt2_3/DFFPOSX1_2/a_34_4# attempt2_3/DFFPOSX1_2/a_22_6# attempt2_3/DFFPOSX1_2/vdd attempt2_3/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1126 attempt2_3/DFFPOSX1_2/a_61_74# attempt2_3/DFFPOSX1_2/a_34_4# attempt2_3/DFFPOSX1_2/vdd attempt2_3/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1127 attempt2_3/DFFPOSX1_2/a_66_6# attempt2_3/DFFPOSX1_2/a_2_6# attempt2_3/DFFPOSX1_2/a_61_74# attempt2_3/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1128 attempt2_3/DFFPOSX1_2/a_76_84# attempt2_3/m1_n35_n168# attempt2_3/DFFPOSX1_2/a_66_6# attempt2_3/DFFPOSX1_2/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1129 attempt2_3/DFFPOSX1_2/vdd attempt2_3/m1_71_n159# attempt2_3/DFFPOSX1_2/a_76_84# attempt2_3/DFFPOSX1_2/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 attempt2_3/DFFPOSX1_2/gnd attempt2_3/m1_n35_n168# attempt2_3/DFFPOSX1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1131 attempt2_3/m1_71_n159# attempt2_3/DFFPOSX1_2/a_66_6# attempt2_3/DFFPOSX1_2/vdd attempt2_3/DFFPOSX1_2/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1132 attempt2_3/DFFPOSX1_2/a_17_6# attempt2_3/m1_n64_n214# attempt2_3/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1133 attempt2_3/DFFPOSX1_2/a_22_6# attempt2_3/DFFPOSX1_2/a_2_6# attempt2_3/DFFPOSX1_2/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1134 attempt2_3/DFFPOSX1_2/a_31_6# attempt2_3/m1_n35_n168# attempt2_3/DFFPOSX1_2/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1135 attempt2_3/DFFPOSX1_2/gnd attempt2_3/DFFPOSX1_2/a_34_4# attempt2_3/DFFPOSX1_2/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1136 attempt2_3/DFFPOSX1_2/a_34_4# attempt2_3/DFFPOSX1_2/a_22_6# attempt2_3/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1137 attempt2_3/DFFPOSX1_2/a_61_6# attempt2_3/DFFPOSX1_2/a_34_4# attempt2_3/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1138 attempt2_3/DFFPOSX1_2/a_66_6# attempt2_3/m1_n35_n168# attempt2_3/DFFPOSX1_2/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1139 attempt2_3/DFFPOSX1_2/a_76_6# attempt2_3/DFFPOSX1_2/a_2_6# attempt2_3/DFFPOSX1_2/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1140 attempt2_3/DFFPOSX1_2/gnd attempt2_3/m1_71_n159# attempt2_3/DFFPOSX1_2/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1141 attempt2_3/m1_71_n159# attempt2_3/DFFPOSX1_2/a_66_6# attempt2_3/DFFPOSX1_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1142 attempt2_3/OR2X1_0/a_9_54# attempt2_3/Input3 attempt2_3/OR2X1_0/a_2_54# attempt2_3/OR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1143 attempt2_3/OR2X1_0/vdd attempt2_3/m1_133_15# attempt2_3/OR2X1_0/a_9_54# attempt2_3/OR2X1_0/vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1144 attempt2_4/Input3 attempt2_3/OR2X1_0/a_2_54# attempt2_3/OR2X1_0/vdd attempt2_3/OR2X1_0/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1145 attempt2_3/OR2X1_0/a_2_54# attempt2_3/Input3 attempt2_3/OR2X1_0/gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=110 ps=62
M1146 attempt2_3/OR2X1_0/gnd attempt2_3/m1_133_15# attempt2_3/OR2X1_0/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 attempt2_4/Input3 attempt2_3/OR2X1_0/a_2_54# attempt2_3/OR2X1_0/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1148 attempt2_3/XOR2X1_0/vdd attempt2_3/m1_n54_n42# attempt2_3/XOR2X1_0/a_2_6# attempt2_3/XOR2X1_0/vdd pfet w=40 l=2
+  ad=560 pd=188 as=200 ps=90
M1149 attempt2_3/XOR2X1_0/a_18_54# attempt2_3/XOR2X1_0/a_13_43# attempt2_3/XOR2X1_0/vdd attempt2_3/XOR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1150 attempt2_3/m1_133_15# attempt2_3/m1_n54_n42# attempt2_3/XOR2X1_0/a_18_54# attempt2_3/XOR2X1_0/vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1151 attempt2_3/XOR2X1_0/a_35_54# attempt2_3/XOR2X1_0/a_2_6# attempt2_3/m1_133_15# attempt2_3/XOR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1152 attempt2_3/XOR2X1_0/vdd attempt2_3/m1_n64_n214# attempt2_3/XOR2X1_0/a_35_54# attempt2_3/XOR2X1_0/vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1153 attempt2_3/XOR2X1_0/a_13_43# attempt2_3/m1_n64_n214# attempt2_3/XOR2X1_0/vdd attempt2_3/XOR2X1_0/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1154 attempt2_3/XOR2X1_0/gnd attempt2_3/m1_n54_n42# attempt2_3/XOR2X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=280 pd=108 as=100 ps=50
M1155 attempt2_3/XOR2X1_0/a_18_6# attempt2_3/XOR2X1_0/a_13_43# attempt2_3/XOR2X1_0/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1156 attempt2_3/m1_133_15# attempt2_3/XOR2X1_0/a_2_6# attempt2_3/XOR2X1_0/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1157 attempt2_3/XOR2X1_0/a_35_6# attempt2_3/m1_n54_n42# attempt2_3/m1_133_15# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1158 attempt2_3/XOR2X1_0/gnd attempt2_3/m1_n64_n214# attempt2_3/XOR2X1_0/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 attempt2_3/XOR2X1_0/a_13_43# attempt2_3/m1_n64_n214# attempt2_3/XOR2X1_0/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1160 attempt2_3/DFFPOSX1_1/vdd attempt2_3/m1_n31_n51# attempt2_3/DFFPOSX1_1/a_2_6# attempt2_3/DFFPOSX1_1/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1161 attempt2_3/DFFPOSX1_1/a_17_74# attempt2_3/m1_n54_n42# attempt2_3/DFFPOSX1_1/vdd attempt2_3/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1162 attempt2_3/DFFPOSX1_1/a_22_6# attempt2_3/m1_n31_n51# attempt2_3/DFFPOSX1_1/a_17_74# attempt2_3/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1163 attempt2_3/DFFPOSX1_1/a_31_74# attempt2_3/DFFPOSX1_1/a_2_6# attempt2_3/DFFPOSX1_1/a_22_6# attempt2_3/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1164 attempt2_3/DFFPOSX1_1/vdd attempt2_3/DFFPOSX1_1/a_34_4# attempt2_3/DFFPOSX1_1/a_31_74# attempt2_3/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1165 attempt2_3/DFFPOSX1_1/a_34_4# attempt2_3/DFFPOSX1_1/a_22_6# attempt2_3/DFFPOSX1_1/vdd attempt2_3/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1166 attempt2_3/DFFPOSX1_1/a_61_74# attempt2_3/DFFPOSX1_1/a_34_4# attempt2_3/DFFPOSX1_1/vdd attempt2_3/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1167 attempt2_3/DFFPOSX1_1/a_66_6# attempt2_3/DFFPOSX1_1/a_2_6# attempt2_3/DFFPOSX1_1/a_61_74# attempt2_3/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1168 attempt2_3/DFFPOSX1_1/a_76_84# attempt2_3/m1_n31_n51# attempt2_3/DFFPOSX1_1/a_66_6# attempt2_3/DFFPOSX1_1/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1169 attempt2_3/DFFPOSX1_1/vdd attempt2_3/m1_n64_n214# attempt2_3/DFFPOSX1_1/a_76_84# attempt2_3/DFFPOSX1_1/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 attempt2_3/DFFPOSX1_1/gnd attempt2_3/m1_n31_n51# attempt2_3/DFFPOSX1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1171 attempt2_3/m1_n64_n214# attempt2_3/DFFPOSX1_1/a_66_6# attempt2_3/DFFPOSX1_1/vdd attempt2_3/DFFPOSX1_1/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1172 attempt2_3/DFFPOSX1_1/a_17_6# attempt2_3/m1_n54_n42# attempt2_3/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1173 attempt2_3/DFFPOSX1_1/a_22_6# attempt2_3/DFFPOSX1_1/a_2_6# attempt2_3/DFFPOSX1_1/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1174 attempt2_3/DFFPOSX1_1/a_31_6# attempt2_3/m1_n31_n51# attempt2_3/DFFPOSX1_1/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1175 attempt2_3/DFFPOSX1_1/gnd attempt2_3/DFFPOSX1_1/a_34_4# attempt2_3/DFFPOSX1_1/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 attempt2_3/DFFPOSX1_1/a_34_4# attempt2_3/DFFPOSX1_1/a_22_6# attempt2_3/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1177 attempt2_3/DFFPOSX1_1/a_61_6# attempt2_3/DFFPOSX1_1/a_34_4# attempt2_3/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1178 attempt2_3/DFFPOSX1_1/a_66_6# attempt2_3/m1_n31_n51# attempt2_3/DFFPOSX1_1/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1179 attempt2_3/DFFPOSX1_1/a_76_6# attempt2_3/DFFPOSX1_1/a_2_6# attempt2_3/DFFPOSX1_1/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1180 attempt2_3/DFFPOSX1_1/gnd attempt2_3/m1_n64_n214# attempt2_3/DFFPOSX1_1/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1181 attempt2_3/m1_n64_n214# attempt2_3/DFFPOSX1_1/a_66_6# attempt2_3/DFFPOSX1_1/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1182 attempt2_3/DFFPOSX1_0/vdd attempt2_3/m1_n29_66# attempt2_3/DFFPOSX1_0/a_2_6# attempt2_3/DFFPOSX1_0/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1183 attempt2_3/DFFPOSX1_0/a_17_74# attempt2_3/Input1 attempt2_3/DFFPOSX1_0/vdd attempt2_3/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1184 attempt2_3/DFFPOSX1_0/a_22_6# attempt2_3/m1_n29_66# attempt2_3/DFFPOSX1_0/a_17_74# attempt2_3/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1185 attempt2_3/DFFPOSX1_0/a_31_74# attempt2_3/DFFPOSX1_0/a_2_6# attempt2_3/DFFPOSX1_0/a_22_6# attempt2_3/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1186 attempt2_3/DFFPOSX1_0/vdd attempt2_3/DFFPOSX1_0/a_34_4# attempt2_3/DFFPOSX1_0/a_31_74# attempt2_3/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 attempt2_3/DFFPOSX1_0/a_34_4# attempt2_3/DFFPOSX1_0/a_22_6# attempt2_3/DFFPOSX1_0/vdd attempt2_3/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1188 attempt2_3/DFFPOSX1_0/a_61_74# attempt2_3/DFFPOSX1_0/a_34_4# attempt2_3/DFFPOSX1_0/vdd attempt2_3/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1189 attempt2_3/DFFPOSX1_0/a_66_6# attempt2_3/DFFPOSX1_0/a_2_6# attempt2_3/DFFPOSX1_0/a_61_74# attempt2_3/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1190 attempt2_3/DFFPOSX1_0/a_76_84# attempt2_3/m1_n29_66# attempt2_3/DFFPOSX1_0/a_66_6# attempt2_3/DFFPOSX1_0/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1191 attempt2_3/DFFPOSX1_0/vdd attempt2_3/m1_n54_n42# attempt2_3/DFFPOSX1_0/a_76_84# attempt2_3/DFFPOSX1_0/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 attempt2_3/DFFPOSX1_0/gnd attempt2_3/m1_n29_66# attempt2_3/DFFPOSX1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1193 attempt2_3/m1_n54_n42# attempt2_3/DFFPOSX1_0/a_66_6# attempt2_3/DFFPOSX1_0/vdd attempt2_3/DFFPOSX1_0/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1194 attempt2_3/DFFPOSX1_0/a_17_6# attempt2_3/Input1 attempt2_3/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1195 attempt2_3/DFFPOSX1_0/a_22_6# attempt2_3/DFFPOSX1_0/a_2_6# attempt2_3/DFFPOSX1_0/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1196 attempt2_3/DFFPOSX1_0/a_31_6# attempt2_3/m1_n29_66# attempt2_3/DFFPOSX1_0/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1197 attempt2_3/DFFPOSX1_0/gnd attempt2_3/DFFPOSX1_0/a_34_4# attempt2_3/DFFPOSX1_0/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 attempt2_3/DFFPOSX1_0/a_34_4# attempt2_3/DFFPOSX1_0/a_22_6# attempt2_3/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1199 attempt2_3/DFFPOSX1_0/a_61_6# attempt2_3/DFFPOSX1_0/a_34_4# attempt2_3/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1200 attempt2_3/DFFPOSX1_0/a_66_6# attempt2_3/m1_n29_66# attempt2_3/DFFPOSX1_0/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1201 attempt2_3/DFFPOSX1_0/a_76_6# attempt2_3/DFFPOSX1_0/a_2_6# attempt2_3/DFFPOSX1_0/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1202 attempt2_3/DFFPOSX1_0/gnd attempt2_3/m1_n54_n42# attempt2_3/DFFPOSX1_0/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1203 attempt2_3/m1_n54_n42# attempt2_3/DFFPOSX1_0/a_66_6# attempt2_3/DFFPOSX1_0/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1204 attempt2_2/OR2X1_1/a_9_54# attempt2_2/m1_133_n102# attempt2_2/OR2X1_1/a_2_54# attempt2_2/OR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1205 attempt2_2/OR2X1_1/vdd attempt2_2/Input2 attempt2_2/OR2X1_1/a_9_54# attempt2_2/OR2X1_1/vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1206 attempt2_3/Input2 attempt2_2/OR2X1_1/a_2_54# attempt2_2/OR2X1_1/vdd attempt2_2/OR2X1_1/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1207 attempt2_2/OR2X1_1/a_2_54# attempt2_2/m1_133_n102# attempt2_2/OR2X1_1/gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=110 ps=62
M1208 attempt2_2/OR2X1_1/gnd attempt2_2/Input2 attempt2_2/OR2X1_1/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 attempt2_3/Input2 attempt2_2/OR2X1_1/a_2_54# attempt2_2/OR2X1_1/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1210 attempt2_2/XOR2X1_1/vdd attempt2_2/m1_n54_n42# attempt2_2/XOR2X1_1/a_2_6# attempt2_2/XOR2X1_1/vdd pfet w=40 l=2
+  ad=560 pd=188 as=200 ps=90
M1211 attempt2_2/XOR2X1_1/a_18_54# attempt2_2/XOR2X1_1/a_13_43# attempt2_2/XOR2X1_1/vdd attempt2_2/XOR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1212 attempt2_2/m1_133_n102# attempt2_2/m1_n54_n42# attempt2_2/XOR2X1_1/a_18_54# attempt2_2/XOR2X1_1/vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1213 attempt2_2/XOR2X1_1/a_35_54# attempt2_2/XOR2X1_1/a_2_6# attempt2_2/m1_133_n102# attempt2_2/XOR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1214 attempt2_2/XOR2X1_1/vdd attempt2_2/m1_71_n159# attempt2_2/XOR2X1_1/a_35_54# attempt2_2/XOR2X1_1/vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 attempt2_2/XOR2X1_1/a_13_43# attempt2_2/m1_71_n159# attempt2_2/XOR2X1_1/vdd attempt2_2/XOR2X1_1/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1216 attempt2_2/XOR2X1_1/gnd attempt2_2/m1_n54_n42# attempt2_2/XOR2X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=280 pd=108 as=100 ps=50
M1217 attempt2_2/XOR2X1_1/a_18_6# attempt2_2/XOR2X1_1/a_13_43# attempt2_2/XOR2X1_1/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1218 attempt2_2/m1_133_n102# attempt2_2/XOR2X1_1/a_2_6# attempt2_2/XOR2X1_1/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1219 attempt2_2/XOR2X1_1/a_35_6# attempt2_2/m1_n54_n42# attempt2_2/m1_133_n102# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1220 attempt2_2/XOR2X1_1/gnd attempt2_2/m1_71_n159# attempt2_2/XOR2X1_1/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1221 attempt2_2/XOR2X1_1/a_13_43# attempt2_2/m1_71_n159# attempt2_2/XOR2X1_1/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1222 attempt2_2/DFFPOSX1_2/vdd attempt2_2/m1_n35_n168# attempt2_2/DFFPOSX1_2/a_2_6# attempt2_2/DFFPOSX1_2/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1223 attempt2_2/DFFPOSX1_2/a_17_74# attempt2_2/m1_n64_n214# attempt2_2/DFFPOSX1_2/vdd attempt2_2/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1224 attempt2_2/DFFPOSX1_2/a_22_6# attempt2_2/m1_n35_n168# attempt2_2/DFFPOSX1_2/a_17_74# attempt2_2/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1225 attempt2_2/DFFPOSX1_2/a_31_74# attempt2_2/DFFPOSX1_2/a_2_6# attempt2_2/DFFPOSX1_2/a_22_6# attempt2_2/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1226 attempt2_2/DFFPOSX1_2/vdd attempt2_2/DFFPOSX1_2/a_34_4# attempt2_2/DFFPOSX1_2/a_31_74# attempt2_2/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 attempt2_2/DFFPOSX1_2/a_34_4# attempt2_2/DFFPOSX1_2/a_22_6# attempt2_2/DFFPOSX1_2/vdd attempt2_2/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1228 attempt2_2/DFFPOSX1_2/a_61_74# attempt2_2/DFFPOSX1_2/a_34_4# attempt2_2/DFFPOSX1_2/vdd attempt2_2/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1229 attempt2_2/DFFPOSX1_2/a_66_6# attempt2_2/DFFPOSX1_2/a_2_6# attempt2_2/DFFPOSX1_2/a_61_74# attempt2_2/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1230 attempt2_2/DFFPOSX1_2/a_76_84# attempt2_2/m1_n35_n168# attempt2_2/DFFPOSX1_2/a_66_6# attempt2_2/DFFPOSX1_2/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1231 attempt2_2/DFFPOSX1_2/vdd attempt2_2/m1_71_n159# attempt2_2/DFFPOSX1_2/a_76_84# attempt2_2/DFFPOSX1_2/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 attempt2_2/DFFPOSX1_2/gnd attempt2_2/m1_n35_n168# attempt2_2/DFFPOSX1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1233 attempt2_2/m1_71_n159# attempt2_2/DFFPOSX1_2/a_66_6# attempt2_2/DFFPOSX1_2/vdd attempt2_2/DFFPOSX1_2/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1234 attempt2_2/DFFPOSX1_2/a_17_6# attempt2_2/m1_n64_n214# attempt2_2/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1235 attempt2_2/DFFPOSX1_2/a_22_6# attempt2_2/DFFPOSX1_2/a_2_6# attempt2_2/DFFPOSX1_2/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1236 attempt2_2/DFFPOSX1_2/a_31_6# attempt2_2/m1_n35_n168# attempt2_2/DFFPOSX1_2/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1237 attempt2_2/DFFPOSX1_2/gnd attempt2_2/DFFPOSX1_2/a_34_4# attempt2_2/DFFPOSX1_2/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1238 attempt2_2/DFFPOSX1_2/a_34_4# attempt2_2/DFFPOSX1_2/a_22_6# attempt2_2/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1239 attempt2_2/DFFPOSX1_2/a_61_6# attempt2_2/DFFPOSX1_2/a_34_4# attempt2_2/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1240 attempt2_2/DFFPOSX1_2/a_66_6# attempt2_2/m1_n35_n168# attempt2_2/DFFPOSX1_2/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1241 attempt2_2/DFFPOSX1_2/a_76_6# attempt2_2/DFFPOSX1_2/a_2_6# attempt2_2/DFFPOSX1_2/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1242 attempt2_2/DFFPOSX1_2/gnd attempt2_2/m1_71_n159# attempt2_2/DFFPOSX1_2/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1243 attempt2_2/m1_71_n159# attempt2_2/DFFPOSX1_2/a_66_6# attempt2_2/DFFPOSX1_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1244 attempt2_2/OR2X1_0/a_9_54# attempt2_2/Input3 attempt2_2/OR2X1_0/a_2_54# attempt2_2/OR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1245 attempt2_2/OR2X1_0/vdd attempt2_2/m1_133_15# attempt2_2/OR2X1_0/a_9_54# attempt2_2/OR2X1_0/vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1246 attempt2_3/Input3 attempt2_2/OR2X1_0/a_2_54# attempt2_2/OR2X1_0/vdd attempt2_2/OR2X1_0/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1247 attempt2_2/OR2X1_0/a_2_54# attempt2_2/Input3 attempt2_2/OR2X1_0/gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=110 ps=62
M1248 attempt2_2/OR2X1_0/gnd attempt2_2/m1_133_15# attempt2_2/OR2X1_0/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1249 attempt2_3/Input3 attempt2_2/OR2X1_0/a_2_54# attempt2_2/OR2X1_0/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1250 attempt2_2/XOR2X1_0/vdd attempt2_2/m1_n54_n42# attempt2_2/XOR2X1_0/a_2_6# attempt2_2/XOR2X1_0/vdd pfet w=40 l=2
+  ad=560 pd=188 as=200 ps=90
M1251 attempt2_2/XOR2X1_0/a_18_54# attempt2_2/XOR2X1_0/a_13_43# attempt2_2/XOR2X1_0/vdd attempt2_2/XOR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1252 attempt2_2/m1_133_15# attempt2_2/m1_n54_n42# attempt2_2/XOR2X1_0/a_18_54# attempt2_2/XOR2X1_0/vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1253 attempt2_2/XOR2X1_0/a_35_54# attempt2_2/XOR2X1_0/a_2_6# attempt2_2/m1_133_15# attempt2_2/XOR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1254 attempt2_2/XOR2X1_0/vdd attempt2_2/m1_n64_n214# attempt2_2/XOR2X1_0/a_35_54# attempt2_2/XOR2X1_0/vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1255 attempt2_2/XOR2X1_0/a_13_43# attempt2_2/m1_n64_n214# attempt2_2/XOR2X1_0/vdd attempt2_2/XOR2X1_0/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1256 attempt2_2/XOR2X1_0/gnd attempt2_2/m1_n54_n42# attempt2_2/XOR2X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=280 pd=108 as=100 ps=50
M1257 attempt2_2/XOR2X1_0/a_18_6# attempt2_2/XOR2X1_0/a_13_43# attempt2_2/XOR2X1_0/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1258 attempt2_2/m1_133_15# attempt2_2/XOR2X1_0/a_2_6# attempt2_2/XOR2X1_0/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1259 attempt2_2/XOR2X1_0/a_35_6# attempt2_2/m1_n54_n42# attempt2_2/m1_133_15# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1260 attempt2_2/XOR2X1_0/gnd attempt2_2/m1_n64_n214# attempt2_2/XOR2X1_0/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1261 attempt2_2/XOR2X1_0/a_13_43# attempt2_2/m1_n64_n214# attempt2_2/XOR2X1_0/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1262 attempt2_2/DFFPOSX1_1/vdd attempt2_2/m1_n31_n51# attempt2_2/DFFPOSX1_1/a_2_6# attempt2_2/DFFPOSX1_1/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1263 attempt2_2/DFFPOSX1_1/a_17_74# attempt2_2/m1_n54_n42# attempt2_2/DFFPOSX1_1/vdd attempt2_2/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1264 attempt2_2/DFFPOSX1_1/a_22_6# attempt2_2/m1_n31_n51# attempt2_2/DFFPOSX1_1/a_17_74# attempt2_2/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1265 attempt2_2/DFFPOSX1_1/a_31_74# attempt2_2/DFFPOSX1_1/a_2_6# attempt2_2/DFFPOSX1_1/a_22_6# attempt2_2/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1266 attempt2_2/DFFPOSX1_1/vdd attempt2_2/DFFPOSX1_1/a_34_4# attempt2_2/DFFPOSX1_1/a_31_74# attempt2_2/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1267 attempt2_2/DFFPOSX1_1/a_34_4# attempt2_2/DFFPOSX1_1/a_22_6# attempt2_2/DFFPOSX1_1/vdd attempt2_2/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1268 attempt2_2/DFFPOSX1_1/a_61_74# attempt2_2/DFFPOSX1_1/a_34_4# attempt2_2/DFFPOSX1_1/vdd attempt2_2/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1269 attempt2_2/DFFPOSX1_1/a_66_6# attempt2_2/DFFPOSX1_1/a_2_6# attempt2_2/DFFPOSX1_1/a_61_74# attempt2_2/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1270 attempt2_2/DFFPOSX1_1/a_76_84# attempt2_2/m1_n31_n51# attempt2_2/DFFPOSX1_1/a_66_6# attempt2_2/DFFPOSX1_1/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1271 attempt2_2/DFFPOSX1_1/vdd attempt2_2/m1_n64_n214# attempt2_2/DFFPOSX1_1/a_76_84# attempt2_2/DFFPOSX1_1/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1272 attempt2_2/DFFPOSX1_1/gnd attempt2_2/m1_n31_n51# attempt2_2/DFFPOSX1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1273 attempt2_2/m1_n64_n214# attempt2_2/DFFPOSX1_1/a_66_6# attempt2_2/DFFPOSX1_1/vdd attempt2_2/DFFPOSX1_1/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1274 attempt2_2/DFFPOSX1_1/a_17_6# attempt2_2/m1_n54_n42# attempt2_2/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1275 attempt2_2/DFFPOSX1_1/a_22_6# attempt2_2/DFFPOSX1_1/a_2_6# attempt2_2/DFFPOSX1_1/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1276 attempt2_2/DFFPOSX1_1/a_31_6# attempt2_2/m1_n31_n51# attempt2_2/DFFPOSX1_1/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1277 attempt2_2/DFFPOSX1_1/gnd attempt2_2/DFFPOSX1_1/a_34_4# attempt2_2/DFFPOSX1_1/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1278 attempt2_2/DFFPOSX1_1/a_34_4# attempt2_2/DFFPOSX1_1/a_22_6# attempt2_2/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1279 attempt2_2/DFFPOSX1_1/a_61_6# attempt2_2/DFFPOSX1_1/a_34_4# attempt2_2/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1280 attempt2_2/DFFPOSX1_1/a_66_6# attempt2_2/m1_n31_n51# attempt2_2/DFFPOSX1_1/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1281 attempt2_2/DFFPOSX1_1/a_76_6# attempt2_2/DFFPOSX1_1/a_2_6# attempt2_2/DFFPOSX1_1/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1282 attempt2_2/DFFPOSX1_1/gnd attempt2_2/m1_n64_n214# attempt2_2/DFFPOSX1_1/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1283 attempt2_2/m1_n64_n214# attempt2_2/DFFPOSX1_1/a_66_6# attempt2_2/DFFPOSX1_1/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1284 attempt2_2/DFFPOSX1_0/vdd attempt2_2/m1_n29_66# attempt2_2/DFFPOSX1_0/a_2_6# attempt2_2/DFFPOSX1_0/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1285 attempt2_2/DFFPOSX1_0/a_17_74# attempt2_2/Input1 attempt2_2/DFFPOSX1_0/vdd attempt2_2/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1286 attempt2_2/DFFPOSX1_0/a_22_6# attempt2_2/m1_n29_66# attempt2_2/DFFPOSX1_0/a_17_74# attempt2_2/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1287 attempt2_2/DFFPOSX1_0/a_31_74# attempt2_2/DFFPOSX1_0/a_2_6# attempt2_2/DFFPOSX1_0/a_22_6# attempt2_2/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1288 attempt2_2/DFFPOSX1_0/vdd attempt2_2/DFFPOSX1_0/a_34_4# attempt2_2/DFFPOSX1_0/a_31_74# attempt2_2/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1289 attempt2_2/DFFPOSX1_0/a_34_4# attempt2_2/DFFPOSX1_0/a_22_6# attempt2_2/DFFPOSX1_0/vdd attempt2_2/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1290 attempt2_2/DFFPOSX1_0/a_61_74# attempt2_2/DFFPOSX1_0/a_34_4# attempt2_2/DFFPOSX1_0/vdd attempt2_2/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1291 attempt2_2/DFFPOSX1_0/a_66_6# attempt2_2/DFFPOSX1_0/a_2_6# attempt2_2/DFFPOSX1_0/a_61_74# attempt2_2/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1292 attempt2_2/DFFPOSX1_0/a_76_84# attempt2_2/m1_n29_66# attempt2_2/DFFPOSX1_0/a_66_6# attempt2_2/DFFPOSX1_0/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1293 attempt2_2/DFFPOSX1_0/vdd attempt2_2/m1_n54_n42# attempt2_2/DFFPOSX1_0/a_76_84# attempt2_2/DFFPOSX1_0/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1294 attempt2_2/DFFPOSX1_0/gnd attempt2_2/m1_n29_66# attempt2_2/DFFPOSX1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1295 attempt2_2/m1_n54_n42# attempt2_2/DFFPOSX1_0/a_66_6# attempt2_2/DFFPOSX1_0/vdd attempt2_2/DFFPOSX1_0/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1296 attempt2_2/DFFPOSX1_0/a_17_6# attempt2_2/Input1 attempt2_2/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1297 attempt2_2/DFFPOSX1_0/a_22_6# attempt2_2/DFFPOSX1_0/a_2_6# attempt2_2/DFFPOSX1_0/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1298 attempt2_2/DFFPOSX1_0/a_31_6# attempt2_2/m1_n29_66# attempt2_2/DFFPOSX1_0/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1299 attempt2_2/DFFPOSX1_0/gnd attempt2_2/DFFPOSX1_0/a_34_4# attempt2_2/DFFPOSX1_0/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1300 attempt2_2/DFFPOSX1_0/a_34_4# attempt2_2/DFFPOSX1_0/a_22_6# attempt2_2/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1301 attempt2_2/DFFPOSX1_0/a_61_6# attempt2_2/DFFPOSX1_0/a_34_4# attempt2_2/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1302 attempt2_2/DFFPOSX1_0/a_66_6# attempt2_2/m1_n29_66# attempt2_2/DFFPOSX1_0/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1303 attempt2_2/DFFPOSX1_0/a_76_6# attempt2_2/DFFPOSX1_0/a_2_6# attempt2_2/DFFPOSX1_0/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1304 attempt2_2/DFFPOSX1_0/gnd attempt2_2/m1_n54_n42# attempt2_2/DFFPOSX1_0/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1305 attempt2_2/m1_n54_n42# attempt2_2/DFFPOSX1_0/a_66_6# attempt2_2/DFFPOSX1_0/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1306 attempt2_1/OR2X1_1/a_9_54# attempt2_1/m1_133_n102# attempt2_1/OR2X1_1/a_2_54# attempt2_1/OR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1307 attempt2_1/OR2X1_1/vdd attempt2_1/Input2 attempt2_1/OR2X1_1/a_9_54# attempt2_1/OR2X1_1/vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1308 attempt2_2/Input2 attempt2_1/OR2X1_1/a_2_54# attempt2_1/OR2X1_1/vdd attempt2_1/OR2X1_1/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1309 attempt2_1/OR2X1_1/a_2_54# attempt2_1/m1_133_n102# attempt2_1/OR2X1_1/gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=110 ps=62
M1310 attempt2_1/OR2X1_1/gnd attempt2_1/Input2 attempt2_1/OR2X1_1/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1311 attempt2_2/Input2 attempt2_1/OR2X1_1/a_2_54# attempt2_1/OR2X1_1/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1312 attempt2_1/XOR2X1_1/vdd attempt2_1/m1_n54_n42# attempt2_1/XOR2X1_1/a_2_6# attempt2_1/XOR2X1_1/vdd pfet w=40 l=2
+  ad=560 pd=188 as=200 ps=90
M1313 attempt2_1/XOR2X1_1/a_18_54# attempt2_1/XOR2X1_1/a_13_43# attempt2_1/XOR2X1_1/vdd attempt2_1/XOR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1314 attempt2_1/m1_133_n102# attempt2_1/m1_n54_n42# attempt2_1/XOR2X1_1/a_18_54# attempt2_1/XOR2X1_1/vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1315 attempt2_1/XOR2X1_1/a_35_54# attempt2_1/XOR2X1_1/a_2_6# attempt2_1/m1_133_n102# attempt2_1/XOR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1316 attempt2_1/XOR2X1_1/vdd attempt2_1/m1_71_n159# attempt2_1/XOR2X1_1/a_35_54# attempt2_1/XOR2X1_1/vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1317 attempt2_1/XOR2X1_1/a_13_43# attempt2_1/m1_71_n159# attempt2_1/XOR2X1_1/vdd attempt2_1/XOR2X1_1/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1318 attempt2_1/XOR2X1_1/gnd attempt2_1/m1_n54_n42# attempt2_1/XOR2X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=280 pd=108 as=100 ps=50
M1319 attempt2_1/XOR2X1_1/a_18_6# attempt2_1/XOR2X1_1/a_13_43# attempt2_1/XOR2X1_1/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1320 attempt2_1/m1_133_n102# attempt2_1/XOR2X1_1/a_2_6# attempt2_1/XOR2X1_1/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1321 attempt2_1/XOR2X1_1/a_35_6# attempt2_1/m1_n54_n42# attempt2_1/m1_133_n102# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1322 attempt2_1/XOR2X1_1/gnd attempt2_1/m1_71_n159# attempt2_1/XOR2X1_1/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1323 attempt2_1/XOR2X1_1/a_13_43# attempt2_1/m1_71_n159# attempt2_1/XOR2X1_1/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1324 attempt2_1/DFFPOSX1_2/vdd attempt2_1/m1_n35_n168# attempt2_1/DFFPOSX1_2/a_2_6# attempt2_1/DFFPOSX1_2/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1325 attempt2_1/DFFPOSX1_2/a_17_74# attempt2_1/m1_n64_n214# attempt2_1/DFFPOSX1_2/vdd attempt2_1/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1326 attempt2_1/DFFPOSX1_2/a_22_6# attempt2_1/m1_n35_n168# attempt2_1/DFFPOSX1_2/a_17_74# attempt2_1/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1327 attempt2_1/DFFPOSX1_2/a_31_74# attempt2_1/DFFPOSX1_2/a_2_6# attempt2_1/DFFPOSX1_2/a_22_6# attempt2_1/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1328 attempt2_1/DFFPOSX1_2/vdd attempt2_1/DFFPOSX1_2/a_34_4# attempt2_1/DFFPOSX1_2/a_31_74# attempt2_1/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1329 attempt2_1/DFFPOSX1_2/a_34_4# attempt2_1/DFFPOSX1_2/a_22_6# attempt2_1/DFFPOSX1_2/vdd attempt2_1/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1330 attempt2_1/DFFPOSX1_2/a_61_74# attempt2_1/DFFPOSX1_2/a_34_4# attempt2_1/DFFPOSX1_2/vdd attempt2_1/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1331 attempt2_1/DFFPOSX1_2/a_66_6# attempt2_1/DFFPOSX1_2/a_2_6# attempt2_1/DFFPOSX1_2/a_61_74# attempt2_1/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1332 attempt2_1/DFFPOSX1_2/a_76_84# attempt2_1/m1_n35_n168# attempt2_1/DFFPOSX1_2/a_66_6# attempt2_1/DFFPOSX1_2/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1333 attempt2_1/DFFPOSX1_2/vdd attempt2_1/m1_71_n159# attempt2_1/DFFPOSX1_2/a_76_84# attempt2_1/DFFPOSX1_2/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1334 attempt2_1/DFFPOSX1_2/gnd attempt2_1/m1_n35_n168# attempt2_1/DFFPOSX1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1335 attempt2_1/m1_71_n159# attempt2_1/DFFPOSX1_2/a_66_6# attempt2_1/DFFPOSX1_2/vdd attempt2_1/DFFPOSX1_2/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1336 attempt2_1/DFFPOSX1_2/a_17_6# attempt2_1/m1_n64_n214# attempt2_1/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1337 attempt2_1/DFFPOSX1_2/a_22_6# attempt2_1/DFFPOSX1_2/a_2_6# attempt2_1/DFFPOSX1_2/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1338 attempt2_1/DFFPOSX1_2/a_31_6# attempt2_1/m1_n35_n168# attempt2_1/DFFPOSX1_2/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1339 attempt2_1/DFFPOSX1_2/gnd attempt2_1/DFFPOSX1_2/a_34_4# attempt2_1/DFFPOSX1_2/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1340 attempt2_1/DFFPOSX1_2/a_34_4# attempt2_1/DFFPOSX1_2/a_22_6# attempt2_1/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1341 attempt2_1/DFFPOSX1_2/a_61_6# attempt2_1/DFFPOSX1_2/a_34_4# attempt2_1/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1342 attempt2_1/DFFPOSX1_2/a_66_6# attempt2_1/m1_n35_n168# attempt2_1/DFFPOSX1_2/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1343 attempt2_1/DFFPOSX1_2/a_76_6# attempt2_1/DFFPOSX1_2/a_2_6# attempt2_1/DFFPOSX1_2/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1344 attempt2_1/DFFPOSX1_2/gnd attempt2_1/m1_71_n159# attempt2_1/DFFPOSX1_2/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1345 attempt2_1/m1_71_n159# attempt2_1/DFFPOSX1_2/a_66_6# attempt2_1/DFFPOSX1_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1346 attempt2_1/OR2X1_0/a_9_54# attempt2_1/Input3 attempt2_1/OR2X1_0/a_2_54# attempt2_1/OR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1347 attempt2_1/OR2X1_0/vdd attempt2_1/m1_133_15# attempt2_1/OR2X1_0/a_9_54# attempt2_1/OR2X1_0/vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1348 attempt2_2/Input3 attempt2_1/OR2X1_0/a_2_54# attempt2_1/OR2X1_0/vdd attempt2_1/OR2X1_0/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1349 attempt2_1/OR2X1_0/a_2_54# attempt2_1/Input3 attempt2_1/OR2X1_0/gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=110 ps=62
M1350 attempt2_1/OR2X1_0/gnd attempt2_1/m1_133_15# attempt2_1/OR2X1_0/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1351 attempt2_2/Input3 attempt2_1/OR2X1_0/a_2_54# attempt2_1/OR2X1_0/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1352 attempt2_1/XOR2X1_0/vdd attempt2_1/m1_n54_n42# attempt2_1/XOR2X1_0/a_2_6# attempt2_1/XOR2X1_0/vdd pfet w=40 l=2
+  ad=560 pd=188 as=200 ps=90
M1353 attempt2_1/XOR2X1_0/a_18_54# attempt2_1/XOR2X1_0/a_13_43# attempt2_1/XOR2X1_0/vdd attempt2_1/XOR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1354 attempt2_1/m1_133_15# attempt2_1/m1_n54_n42# attempt2_1/XOR2X1_0/a_18_54# attempt2_1/XOR2X1_0/vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1355 attempt2_1/XOR2X1_0/a_35_54# attempt2_1/XOR2X1_0/a_2_6# attempt2_1/m1_133_15# attempt2_1/XOR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1356 attempt2_1/XOR2X1_0/vdd attempt2_1/m1_n64_n214# attempt2_1/XOR2X1_0/a_35_54# attempt2_1/XOR2X1_0/vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1357 attempt2_1/XOR2X1_0/a_13_43# attempt2_1/m1_n64_n214# attempt2_1/XOR2X1_0/vdd attempt2_1/XOR2X1_0/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1358 attempt2_1/XOR2X1_0/gnd attempt2_1/m1_n54_n42# attempt2_1/XOR2X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=280 pd=108 as=100 ps=50
M1359 attempt2_1/XOR2X1_0/a_18_6# attempt2_1/XOR2X1_0/a_13_43# attempt2_1/XOR2X1_0/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1360 attempt2_1/m1_133_15# attempt2_1/XOR2X1_0/a_2_6# attempt2_1/XOR2X1_0/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1361 attempt2_1/XOR2X1_0/a_35_6# attempt2_1/m1_n54_n42# attempt2_1/m1_133_15# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1362 attempt2_1/XOR2X1_0/gnd attempt2_1/m1_n64_n214# attempt2_1/XOR2X1_0/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1363 attempt2_1/XOR2X1_0/a_13_43# attempt2_1/m1_n64_n214# attempt2_1/XOR2X1_0/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1364 attempt2_1/DFFPOSX1_1/vdd attempt2_1/m1_n31_n51# attempt2_1/DFFPOSX1_1/a_2_6# attempt2_1/DFFPOSX1_1/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1365 attempt2_1/DFFPOSX1_1/a_17_74# attempt2_1/m1_n54_n42# attempt2_1/DFFPOSX1_1/vdd attempt2_1/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1366 attempt2_1/DFFPOSX1_1/a_22_6# attempt2_1/m1_n31_n51# attempt2_1/DFFPOSX1_1/a_17_74# attempt2_1/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1367 attempt2_1/DFFPOSX1_1/a_31_74# attempt2_1/DFFPOSX1_1/a_2_6# attempt2_1/DFFPOSX1_1/a_22_6# attempt2_1/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1368 attempt2_1/DFFPOSX1_1/vdd attempt2_1/DFFPOSX1_1/a_34_4# attempt2_1/DFFPOSX1_1/a_31_74# attempt2_1/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1369 attempt2_1/DFFPOSX1_1/a_34_4# attempt2_1/DFFPOSX1_1/a_22_6# attempt2_1/DFFPOSX1_1/vdd attempt2_1/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1370 attempt2_1/DFFPOSX1_1/a_61_74# attempt2_1/DFFPOSX1_1/a_34_4# attempt2_1/DFFPOSX1_1/vdd attempt2_1/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1371 attempt2_1/DFFPOSX1_1/a_66_6# attempt2_1/DFFPOSX1_1/a_2_6# attempt2_1/DFFPOSX1_1/a_61_74# attempt2_1/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1372 attempt2_1/DFFPOSX1_1/a_76_84# attempt2_1/m1_n31_n51# attempt2_1/DFFPOSX1_1/a_66_6# attempt2_1/DFFPOSX1_1/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1373 attempt2_1/DFFPOSX1_1/vdd attempt2_1/m1_n64_n214# attempt2_1/DFFPOSX1_1/a_76_84# attempt2_1/DFFPOSX1_1/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1374 attempt2_1/DFFPOSX1_1/gnd attempt2_1/m1_n31_n51# attempt2_1/DFFPOSX1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1375 attempt2_1/m1_n64_n214# attempt2_1/DFFPOSX1_1/a_66_6# attempt2_1/DFFPOSX1_1/vdd attempt2_1/DFFPOSX1_1/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1376 attempt2_1/DFFPOSX1_1/a_17_6# attempt2_1/m1_n54_n42# attempt2_1/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1377 attempt2_1/DFFPOSX1_1/a_22_6# attempt2_1/DFFPOSX1_1/a_2_6# attempt2_1/DFFPOSX1_1/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1378 attempt2_1/DFFPOSX1_1/a_31_6# attempt2_1/m1_n31_n51# attempt2_1/DFFPOSX1_1/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1379 attempt2_1/DFFPOSX1_1/gnd attempt2_1/DFFPOSX1_1/a_34_4# attempt2_1/DFFPOSX1_1/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1380 attempt2_1/DFFPOSX1_1/a_34_4# attempt2_1/DFFPOSX1_1/a_22_6# attempt2_1/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1381 attempt2_1/DFFPOSX1_1/a_61_6# attempt2_1/DFFPOSX1_1/a_34_4# attempt2_1/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1382 attempt2_1/DFFPOSX1_1/a_66_6# attempt2_1/m1_n31_n51# attempt2_1/DFFPOSX1_1/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1383 attempt2_1/DFFPOSX1_1/a_76_6# attempt2_1/DFFPOSX1_1/a_2_6# attempt2_1/DFFPOSX1_1/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1384 attempt2_1/DFFPOSX1_1/gnd attempt2_1/m1_n64_n214# attempt2_1/DFFPOSX1_1/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1385 attempt2_1/m1_n64_n214# attempt2_1/DFFPOSX1_1/a_66_6# attempt2_1/DFFPOSX1_1/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1386 attempt2_1/DFFPOSX1_0/vdd attempt2_1/m1_n29_66# attempt2_1/DFFPOSX1_0/a_2_6# attempt2_1/DFFPOSX1_0/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1387 attempt2_1/DFFPOSX1_0/a_17_74# attempt2_1/Input1 attempt2_1/DFFPOSX1_0/vdd attempt2_1/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1388 attempt2_1/DFFPOSX1_0/a_22_6# attempt2_1/m1_n29_66# attempt2_1/DFFPOSX1_0/a_17_74# attempt2_1/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1389 attempt2_1/DFFPOSX1_0/a_31_74# attempt2_1/DFFPOSX1_0/a_2_6# attempt2_1/DFFPOSX1_0/a_22_6# attempt2_1/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1390 attempt2_1/DFFPOSX1_0/vdd attempt2_1/DFFPOSX1_0/a_34_4# attempt2_1/DFFPOSX1_0/a_31_74# attempt2_1/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1391 attempt2_1/DFFPOSX1_0/a_34_4# attempt2_1/DFFPOSX1_0/a_22_6# attempt2_1/DFFPOSX1_0/vdd attempt2_1/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1392 attempt2_1/DFFPOSX1_0/a_61_74# attempt2_1/DFFPOSX1_0/a_34_4# attempt2_1/DFFPOSX1_0/vdd attempt2_1/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1393 attempt2_1/DFFPOSX1_0/a_66_6# attempt2_1/DFFPOSX1_0/a_2_6# attempt2_1/DFFPOSX1_0/a_61_74# attempt2_1/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1394 attempt2_1/DFFPOSX1_0/a_76_84# attempt2_1/m1_n29_66# attempt2_1/DFFPOSX1_0/a_66_6# attempt2_1/DFFPOSX1_0/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1395 attempt2_1/DFFPOSX1_0/vdd attempt2_1/m1_n54_n42# attempt2_1/DFFPOSX1_0/a_76_84# attempt2_1/DFFPOSX1_0/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1396 attempt2_1/DFFPOSX1_0/gnd attempt2_1/m1_n29_66# attempt2_1/DFFPOSX1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1397 attempt2_1/m1_n54_n42# attempt2_1/DFFPOSX1_0/a_66_6# attempt2_1/DFFPOSX1_0/vdd attempt2_1/DFFPOSX1_0/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1398 attempt2_1/DFFPOSX1_0/a_17_6# attempt2_1/Input1 attempt2_1/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1399 attempt2_1/DFFPOSX1_0/a_22_6# attempt2_1/DFFPOSX1_0/a_2_6# attempt2_1/DFFPOSX1_0/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1400 attempt2_1/DFFPOSX1_0/a_31_6# attempt2_1/m1_n29_66# attempt2_1/DFFPOSX1_0/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1401 attempt2_1/DFFPOSX1_0/gnd attempt2_1/DFFPOSX1_0/a_34_4# attempt2_1/DFFPOSX1_0/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1402 attempt2_1/DFFPOSX1_0/a_34_4# attempt2_1/DFFPOSX1_0/a_22_6# attempt2_1/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1403 attempt2_1/DFFPOSX1_0/a_61_6# attempt2_1/DFFPOSX1_0/a_34_4# attempt2_1/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1404 attempt2_1/DFFPOSX1_0/a_66_6# attempt2_1/m1_n29_66# attempt2_1/DFFPOSX1_0/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1405 attempt2_1/DFFPOSX1_0/a_76_6# attempt2_1/DFFPOSX1_0/a_2_6# attempt2_1/DFFPOSX1_0/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1406 attempt2_1/DFFPOSX1_0/gnd attempt2_1/m1_n54_n42# attempt2_1/DFFPOSX1_0/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1407 attempt2_1/m1_n54_n42# attempt2_1/DFFPOSX1_0/a_66_6# attempt2_1/DFFPOSX1_0/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1408 attempt2_0/OR2X1_1/a_9_54# attempt2_0/m1_133_n102# attempt2_0/OR2X1_1/a_2_54# attempt2_0/OR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1409 attempt2_0/OR2X1_1/vdd attempt2_0/Input2 attempt2_0/OR2X1_1/a_9_54# attempt2_0/OR2X1_1/vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1410 attempt2_1/Input2 attempt2_0/OR2X1_1/a_2_54# attempt2_0/OR2X1_1/vdd attempt2_0/OR2X1_1/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1411 attempt2_0/OR2X1_1/a_2_54# attempt2_0/m1_133_n102# attempt2_0/OR2X1_1/gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=110 ps=62
M1412 attempt2_0/OR2X1_1/gnd attempt2_0/Input2 attempt2_0/OR2X1_1/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1413 attempt2_1/Input2 attempt2_0/OR2X1_1/a_2_54# attempt2_0/OR2X1_1/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1414 attempt2_0/XOR2X1_1/vdd attempt2_0/m1_n54_n42# attempt2_0/XOR2X1_1/a_2_6# attempt2_0/XOR2X1_1/vdd pfet w=40 l=2
+  ad=560 pd=188 as=200 ps=90
M1415 attempt2_0/XOR2X1_1/a_18_54# attempt2_0/XOR2X1_1/a_13_43# attempt2_0/XOR2X1_1/vdd attempt2_0/XOR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1416 attempt2_0/m1_133_n102# attempt2_0/m1_n54_n42# attempt2_0/XOR2X1_1/a_18_54# attempt2_0/XOR2X1_1/vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1417 attempt2_0/XOR2X1_1/a_35_54# attempt2_0/XOR2X1_1/a_2_6# attempt2_0/m1_133_n102# attempt2_0/XOR2X1_1/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1418 attempt2_0/XOR2X1_1/vdd attempt2_0/m1_71_n159# attempt2_0/XOR2X1_1/a_35_54# attempt2_0/XOR2X1_1/vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1419 attempt2_0/XOR2X1_1/a_13_43# attempt2_0/m1_71_n159# attempt2_0/XOR2X1_1/vdd attempt2_0/XOR2X1_1/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1420 attempt2_0/XOR2X1_1/gnd attempt2_0/m1_n54_n42# attempt2_0/XOR2X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=280 pd=108 as=100 ps=50
M1421 attempt2_0/XOR2X1_1/a_18_6# attempt2_0/XOR2X1_1/a_13_43# attempt2_0/XOR2X1_1/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1422 attempt2_0/m1_133_n102# attempt2_0/XOR2X1_1/a_2_6# attempt2_0/XOR2X1_1/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1423 attempt2_0/XOR2X1_1/a_35_6# attempt2_0/m1_n54_n42# attempt2_0/m1_133_n102# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1424 attempt2_0/XOR2X1_1/gnd attempt2_0/m1_71_n159# attempt2_0/XOR2X1_1/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1425 attempt2_0/XOR2X1_1/a_13_43# attempt2_0/m1_71_n159# attempt2_0/XOR2X1_1/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1426 attempt2_0/DFFPOSX1_2/vdd attempt2_0/m1_n35_n168# attempt2_0/DFFPOSX1_2/a_2_6# attempt2_0/DFFPOSX1_2/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1427 attempt2_0/DFFPOSX1_2/a_17_74# attempt2_0/m1_n64_n214# attempt2_0/DFFPOSX1_2/vdd attempt2_0/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1428 attempt2_0/DFFPOSX1_2/a_22_6# attempt2_0/m1_n35_n168# attempt2_0/DFFPOSX1_2/a_17_74# attempt2_0/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1429 attempt2_0/DFFPOSX1_2/a_31_74# attempt2_0/DFFPOSX1_2/a_2_6# attempt2_0/DFFPOSX1_2/a_22_6# attempt2_0/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1430 attempt2_0/DFFPOSX1_2/vdd attempt2_0/DFFPOSX1_2/a_34_4# attempt2_0/DFFPOSX1_2/a_31_74# attempt2_0/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1431 attempt2_0/DFFPOSX1_2/a_34_4# attempt2_0/DFFPOSX1_2/a_22_6# attempt2_0/DFFPOSX1_2/vdd attempt2_0/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1432 attempt2_0/DFFPOSX1_2/a_61_74# attempt2_0/DFFPOSX1_2/a_34_4# attempt2_0/DFFPOSX1_2/vdd attempt2_0/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1433 attempt2_0/DFFPOSX1_2/a_66_6# attempt2_0/DFFPOSX1_2/a_2_6# attempt2_0/DFFPOSX1_2/a_61_74# attempt2_0/DFFPOSX1_2/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1434 attempt2_0/DFFPOSX1_2/a_76_84# attempt2_0/m1_n35_n168# attempt2_0/DFFPOSX1_2/a_66_6# attempt2_0/DFFPOSX1_2/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1435 attempt2_0/DFFPOSX1_2/vdd attempt2_0/m1_71_n159# attempt2_0/DFFPOSX1_2/a_76_84# attempt2_0/DFFPOSX1_2/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1436 attempt2_0/DFFPOSX1_2/gnd attempt2_0/m1_n35_n168# attempt2_0/DFFPOSX1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1437 attempt2_0/m1_71_n159# attempt2_0/DFFPOSX1_2/a_66_6# attempt2_0/DFFPOSX1_2/vdd attempt2_0/DFFPOSX1_2/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1438 attempt2_0/DFFPOSX1_2/a_17_6# attempt2_0/m1_n64_n214# attempt2_0/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1439 attempt2_0/DFFPOSX1_2/a_22_6# attempt2_0/DFFPOSX1_2/a_2_6# attempt2_0/DFFPOSX1_2/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1440 attempt2_0/DFFPOSX1_2/a_31_6# attempt2_0/m1_n35_n168# attempt2_0/DFFPOSX1_2/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1441 attempt2_0/DFFPOSX1_2/gnd attempt2_0/DFFPOSX1_2/a_34_4# attempt2_0/DFFPOSX1_2/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1442 attempt2_0/DFFPOSX1_2/a_34_4# attempt2_0/DFFPOSX1_2/a_22_6# attempt2_0/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1443 attempt2_0/DFFPOSX1_2/a_61_6# attempt2_0/DFFPOSX1_2/a_34_4# attempt2_0/DFFPOSX1_2/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1444 attempt2_0/DFFPOSX1_2/a_66_6# attempt2_0/m1_n35_n168# attempt2_0/DFFPOSX1_2/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1445 attempt2_0/DFFPOSX1_2/a_76_6# attempt2_0/DFFPOSX1_2/a_2_6# attempt2_0/DFFPOSX1_2/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1446 attempt2_0/DFFPOSX1_2/gnd attempt2_0/m1_71_n159# attempt2_0/DFFPOSX1_2/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1447 attempt2_0/m1_71_n159# attempt2_0/DFFPOSX1_2/a_66_6# attempt2_0/DFFPOSX1_2/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1448 attempt2_0/OR2X1_0/a_9_54# attempt2_0/Input3 attempt2_0/OR2X1_0/a_2_54# attempt2_0/OR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=200 ps=90
M1449 attempt2_0/OR2X1_0/vdd attempt2_0/m1_133_15# attempt2_0/OR2X1_0/a_9_54# attempt2_0/OR2X1_0/vdd pfet w=40 l=2
+  ad=220 pd=92 as=0 ps=0
M1450 attempt2_1/Input3 attempt2_0/OR2X1_0/a_2_54# attempt2_0/OR2X1_0/vdd attempt2_0/OR2X1_0/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1451 attempt2_0/OR2X1_0/a_2_54# attempt2_0/Input3 attempt2_0/OR2X1_0/gnd Gnd nfet w=10 l=2
+  ad=60 pd=32 as=110 ps=62
M1452 attempt2_0/OR2X1_0/gnd attempt2_0/m1_133_15# attempt2_0/OR2X1_0/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1453 attempt2_1/Input3 attempt2_0/OR2X1_0/a_2_54# attempt2_0/OR2X1_0/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1454 attempt2_0/XOR2X1_0/vdd attempt2_0/m1_n54_n42# attempt2_0/XOR2X1_0/a_2_6# attempt2_0/XOR2X1_0/vdd pfet w=40 l=2
+  ad=560 pd=188 as=200 ps=90
M1455 attempt2_0/XOR2X1_0/a_18_54# attempt2_0/XOR2X1_0/a_13_43# attempt2_0/XOR2X1_0/vdd attempt2_0/XOR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1456 attempt2_0/m1_133_15# attempt2_0/m1_n54_n42# attempt2_0/XOR2X1_0/a_18_54# attempt2_0/XOR2X1_0/vdd pfet w=40 l=2
+  ad=400 pd=100 as=0 ps=0
M1457 attempt2_0/XOR2X1_0/a_35_54# attempt2_0/XOR2X1_0/a_2_6# attempt2_0/m1_133_15# attempt2_0/XOR2X1_0/vdd pfet w=40 l=2
+  ad=120 pd=86 as=0 ps=0
M1458 attempt2_0/XOR2X1_0/vdd attempt2_0/m1_n64_n214# attempt2_0/XOR2X1_0/a_35_54# attempt2_0/XOR2X1_0/vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1459 attempt2_0/XOR2X1_0/a_13_43# attempt2_0/m1_n64_n214# attempt2_0/XOR2X1_0/vdd attempt2_0/XOR2X1_0/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1460 attempt2_0/XOR2X1_0/gnd attempt2_0/m1_n54_n42# attempt2_0/XOR2X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=280 pd=108 as=100 ps=50
M1461 attempt2_0/XOR2X1_0/a_18_6# attempt2_0/XOR2X1_0/a_13_43# attempt2_0/XOR2X1_0/gnd Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1462 attempt2_0/m1_133_15# attempt2_0/XOR2X1_0/a_2_6# attempt2_0/XOR2X1_0/a_18_6# Gnd nfet w=20 l=2
+  ad=200 pd=60 as=0 ps=0
M1463 attempt2_0/XOR2X1_0/a_35_6# attempt2_0/m1_n54_n42# attempt2_0/m1_133_15# Gnd nfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1464 attempt2_0/XOR2X1_0/gnd attempt2_0/m1_n64_n214# attempt2_0/XOR2X1_0/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1465 attempt2_0/XOR2X1_0/a_13_43# attempt2_0/m1_n64_n214# attempt2_0/XOR2X1_0/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1466 attempt2_0/DFFPOSX1_1/vdd attempt2_0/m1_n31_n51# attempt2_0/DFFPOSX1_1/a_2_6# attempt2_0/DFFPOSX1_1/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1467 attempt2_0/DFFPOSX1_1/a_17_74# attempt2_0/m1_n54_n42# attempt2_0/DFFPOSX1_1/vdd attempt2_0/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1468 attempt2_0/DFFPOSX1_1/a_22_6# attempt2_0/m1_n31_n51# attempt2_0/DFFPOSX1_1/a_17_74# attempt2_0/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1469 attempt2_0/DFFPOSX1_1/a_31_74# attempt2_0/DFFPOSX1_1/a_2_6# attempt2_0/DFFPOSX1_1/a_22_6# attempt2_0/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1470 attempt2_0/DFFPOSX1_1/vdd attempt2_0/DFFPOSX1_1/a_34_4# attempt2_0/DFFPOSX1_1/a_31_74# attempt2_0/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1471 attempt2_0/DFFPOSX1_1/a_34_4# attempt2_0/DFFPOSX1_1/a_22_6# attempt2_0/DFFPOSX1_1/vdd attempt2_0/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1472 attempt2_0/DFFPOSX1_1/a_61_74# attempt2_0/DFFPOSX1_1/a_34_4# attempt2_0/DFFPOSX1_1/vdd attempt2_0/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1473 attempt2_0/DFFPOSX1_1/a_66_6# attempt2_0/DFFPOSX1_1/a_2_6# attempt2_0/DFFPOSX1_1/a_61_74# attempt2_0/DFFPOSX1_1/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1474 attempt2_0/DFFPOSX1_1/a_76_84# attempt2_0/m1_n31_n51# attempt2_0/DFFPOSX1_1/a_66_6# attempt2_0/DFFPOSX1_1/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1475 attempt2_0/DFFPOSX1_1/vdd attempt2_0/m1_n64_n214# attempt2_0/DFFPOSX1_1/a_76_84# attempt2_0/DFFPOSX1_1/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1476 attempt2_0/DFFPOSX1_1/gnd attempt2_0/m1_n31_n51# attempt2_0/DFFPOSX1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1477 attempt2_0/m1_n64_n214# attempt2_0/DFFPOSX1_1/a_66_6# attempt2_0/DFFPOSX1_1/vdd attempt2_0/DFFPOSX1_1/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1478 attempt2_0/DFFPOSX1_1/a_17_6# attempt2_0/m1_n54_n42# attempt2_0/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1479 attempt2_0/DFFPOSX1_1/a_22_6# attempt2_0/DFFPOSX1_1/a_2_6# attempt2_0/DFFPOSX1_1/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1480 attempt2_0/DFFPOSX1_1/a_31_6# attempt2_0/m1_n31_n51# attempt2_0/DFFPOSX1_1/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1481 attempt2_0/DFFPOSX1_1/gnd attempt2_0/DFFPOSX1_1/a_34_4# attempt2_0/DFFPOSX1_1/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1482 attempt2_0/DFFPOSX1_1/a_34_4# attempt2_0/DFFPOSX1_1/a_22_6# attempt2_0/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1483 attempt2_0/DFFPOSX1_1/a_61_6# attempt2_0/DFFPOSX1_1/a_34_4# attempt2_0/DFFPOSX1_1/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1484 attempt2_0/DFFPOSX1_1/a_66_6# attempt2_0/m1_n31_n51# attempt2_0/DFFPOSX1_1/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1485 attempt2_0/DFFPOSX1_1/a_76_6# attempt2_0/DFFPOSX1_1/a_2_6# attempt2_0/DFFPOSX1_1/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1486 attempt2_0/DFFPOSX1_1/gnd attempt2_0/m1_n64_n214# attempt2_0/DFFPOSX1_1/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1487 attempt2_0/m1_n64_n214# attempt2_0/DFFPOSX1_1/a_66_6# attempt2_0/DFFPOSX1_1/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1488 attempt2_0/DFFPOSX1_0/vdd attempt2_0/m1_n29_66# attempt2_0/DFFPOSX1_0/a_2_6# attempt2_0/DFFPOSX1_0/vdd pfet w=40 l=2
+  ad=650 pd=286 as=200 ps=90
M1489 attempt2_0/DFFPOSX1_0/a_17_74# attempt2_0/Input1 attempt2_0/DFFPOSX1_0/vdd attempt2_0/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1490 attempt2_0/DFFPOSX1_0/a_22_6# attempt2_0/m1_n29_66# attempt2_0/DFFPOSX1_0/a_17_74# attempt2_0/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1491 attempt2_0/DFFPOSX1_0/a_31_74# attempt2_0/DFFPOSX1_0/a_2_6# attempt2_0/DFFPOSX1_0/a_22_6# attempt2_0/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=80 pd=48 as=0 ps=0
M1492 attempt2_0/DFFPOSX1_0/vdd attempt2_0/DFFPOSX1_0/a_34_4# attempt2_0/DFFPOSX1_0/a_31_74# attempt2_0/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1493 attempt2_0/DFFPOSX1_0/a_34_4# attempt2_0/DFFPOSX1_0/a_22_6# attempt2_0/DFFPOSX1_0/vdd attempt2_0/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1494 attempt2_0/DFFPOSX1_0/a_61_74# attempt2_0/DFFPOSX1_0/a_34_4# attempt2_0/DFFPOSX1_0/vdd attempt2_0/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=60 pd=46 as=0 ps=0
M1495 attempt2_0/DFFPOSX1_0/a_66_6# attempt2_0/DFFPOSX1_0/a_2_6# attempt2_0/DFFPOSX1_0/a_61_74# attempt2_0/DFFPOSX1_0/vdd pfet w=20 l=2
+  ad=150 pd=56 as=0 ps=0
M1496 attempt2_0/DFFPOSX1_0/a_76_84# attempt2_0/m1_n29_66# attempt2_0/DFFPOSX1_0/a_66_6# attempt2_0/DFFPOSX1_0/vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1497 attempt2_0/DFFPOSX1_0/vdd attempt2_0/m1_n54_n42# attempt2_0/DFFPOSX1_0/a_76_84# attempt2_0/DFFPOSX1_0/vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1498 attempt2_0/DFFPOSX1_0/gnd attempt2_0/m1_n29_66# attempt2_0/DFFPOSX1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=340 pd=168 as=100 ps=50
M1499 attempt2_0/m1_n54_n42# attempt2_0/DFFPOSX1_0/a_66_6# attempt2_0/DFFPOSX1_0/vdd attempt2_0/DFFPOSX1_0/vdd pfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1500 attempt2_0/DFFPOSX1_0/a_17_6# attempt2_0/Input1 attempt2_0/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1501 attempt2_0/DFFPOSX1_0/a_22_6# attempt2_0/DFFPOSX1_0/a_2_6# attempt2_0/DFFPOSX1_0/a_17_6# Gnd nfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1502 attempt2_0/DFFPOSX1_0/a_31_6# attempt2_0/m1_n29_66# attempt2_0/DFFPOSX1_0/a_22_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1503 attempt2_0/DFFPOSX1_0/gnd attempt2_0/DFFPOSX1_0/a_34_4# attempt2_0/DFFPOSX1_0/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1504 attempt2_0/DFFPOSX1_0/a_34_4# attempt2_0/DFFPOSX1_0/a_22_6# attempt2_0/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1505 attempt2_0/DFFPOSX1_0/a_61_6# attempt2_0/DFFPOSX1_0/a_34_4# attempt2_0/DFFPOSX1_0/gnd Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1506 attempt2_0/DFFPOSX1_0/a_66_6# attempt2_0/m1_n29_66# attempt2_0/DFFPOSX1_0/a_61_6# Gnd nfet w=10 l=2
+  ad=80 pd=36 as=0 ps=0
M1507 attempt2_0/DFFPOSX1_0/a_76_6# attempt2_0/DFFPOSX1_0/a_2_6# attempt2_0/DFFPOSX1_0/a_66_6# Gnd nfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1508 attempt2_0/DFFPOSX1_0/gnd attempt2_0/m1_n54_n42# attempt2_0/DFFPOSX1_0/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1509 attempt2_0/m1_n54_n42# attempt2_0/DFFPOSX1_0/a_66_6# attempt2_0/DFFPOSX1_0/gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 attempt2_2/DFFPOSX1_2/vdd attempt2_2/DFFPOSX1_2/a_2_6# 4.88fF
C1 attempt2_4/DFFPOSX1_2/a_2_6# attempt2_4/DFFPOSX1_2/vdd 4.88fF
C2 attempt2_1/m1_n64_n214# attempt2_1/DFFPOSX1_1/vdd 2.20fF
C3 attempt2_0/DFFPOSX1_2/vdd attempt2_0/DFFPOSX1_2/a_34_4# 2.48fF
C4 attempt2_4/OR2X1_1/a_2_54# attempt2_4/OR2X1_1/vdd 2.08fF
C5 attempt2_2/DFFPOSX1_1/vdd attempt2_2/DFFPOSX1_1/a_22_6# 2.40fF
C6 attempt2_4/m1_n64_n214# attempt2_4/DFFPOSX1_1/vdd 2.20fF
C7 attempt2_1/DFFPOSX1_0/vdd attempt2_1/DFFPOSX1_0/a_2_6# 4.88fF
C8 attempt2_3/DFFPOSX1_2/vdd attempt2_3/DFFPOSX1_2/a_2_6# 4.88fF
C9 attempt2_2/DFFPOSX1_2/vdd attempt2_2/DFFPOSX1_2/a_34_4# 2.48fF
C10 attempt2_0/DFFPOSX1_0/vdd attempt2_0/m1_n29_66# 2.41fF
C11 attempt2_4/DFFPOSX1_0/vdd attempt2_4/m1_n29_66# 2.41fF
C12 attempt2_1/DFFPOSX1_2/vdd attempt2_1/m1_n35_n168# 2.41fF
C13 attempt2_3/DFFPOSX1_1/vdd attempt2_3/DFFPOSX1_1/a_2_6# 4.88fF
C14 attempt2_4/DFFPOSX1_1/vdd attempt2_4/m1_n31_n51# 2.41fF
C15 attempt2_2/DFFPOSX1_0/vdd attempt2_2/m1_n29_66# 2.41fF
C16 attempt2_1/DFFPOSX1_0/vdd attempt2_1/DFFPOSX1_0/a_34_4# 2.48fF
C17 attempt2_1/DFFPOSX1_1/vdd attempt2_1/DFFPOSX1_1/a_2_6# 4.88fF
C18 attempt2_4/m1_n35_n168# attempt2_4/DFFPOSX1_2/vdd 2.41fF
C19 attempt2_2/DFFPOSX1_0/vdd attempt2_2/DFFPOSX1_0/a_22_6# 2.40fF
C20 attempt2_1/OR2X1_0/vdd attempt2_1/OR2X1_0/a_2_54# 2.08fF
C21 attempt2_0/DFFPOSX1_2/vdd attempt2_0/DFFPOSX1_2/a_22_6# 2.40fF
C22 attempt2_1/OR2X1_1/vdd attempt2_1/OR2X1_1/a_2_54# 2.08fF
C23 attempt2_2/DFFPOSX1_2/vdd attempt2_2/DFFPOSX1_2/a_22_6# 2.40fF
C24 attempt2_4/DFFPOSX1_0/vdd attempt2_4/DFFPOSX1_0/a_2_6# 4.88fF
C25 attempt2_0/DFFPOSX1_1/vdd attempt2_0/m1_n31_n51# 2.41fF
C26 attempt2_0/m1_71_n159# attempt2_0/DFFPOSX1_2/vdd 2.20fF
C27 attempt2_3/DFFPOSX1_1/vdd attempt2_3/DFFPOSX1_1/a_34_4# 2.48fF
C28 attempt2_4/DFFPOSX1_1/vdd attempt2_4/DFFPOSX1_1/a_2_6# 4.88fF
C29 attempt2_2/DFFPOSX1_1/vdd attempt2_2/m1_n31_n51# 2.41fF
C30 attempt2_1/DFFPOSX1_0/vdd attempt2_1/DFFPOSX1_0/a_22_6# 2.40fF
C31 attempt2_1/DFFPOSX1_1/vdd attempt2_1/DFFPOSX1_1/a_34_4# 2.48fF
C32 attempt2_2/m1_71_n159# attempt2_2/DFFPOSX1_2/vdd 2.20fF
C33 attempt2_3/DFFPOSX1_0/vdd attempt2_3/DFFPOSX1_0/a_2_6# 4.88fF
C34 attempt2_0/DFFPOSX1_0/vdd attempt2_0/DFFPOSX1_0/a_2_6# 4.88fF
C35 attempt2_3/m1_71_n159# attempt2_3/DFFPOSX1_2/vdd 2.20fF
C36 attempt2_4/DFFPOSX1_0/vdd attempt2_4/DFFPOSX1_0/a_34_4# 2.48fF
C37 attempt2_2/m1_n54_n42# attempt2_2/DFFPOSX1_0/vdd 2.20fF
C38 attempt2_4/DFFPOSX1_1/vdd attempt2_4/DFFPOSX1_1/a_34_4# 2.48fF
C39 attempt2_3/OR2X1_0/vdd attempt2_3/OR2X1_0/a_2_54# 2.08fF
C40 attempt2_4/DFFPOSX1_0/vdd attempt2_4/DFFPOSX1_0/a_22_6# 2.40fF
C41 attempt2_2/m1_n64_n214# attempt2_2/DFFPOSX1_1/vdd 2.20fF
C42 attempt2_3/DFFPOSX1_2/a_34_4# attempt2_3/DFFPOSX1_2/vdd 2.48fF
C43 attempt2_1/DFFPOSX1_2/vdd attempt2_1/DFFPOSX1_2/a_2_6# 4.88fF
C44 attempt2_1/m1_n54_n42# attempt2_1/DFFPOSX1_0/vdd 2.20fF
C45 attempt2_0/DFFPOSX1_2/vdd attempt2_0/m1_n35_n168# 2.41fF
C46 attempt2_3/DFFPOSX1_1/vdd attempt2_3/DFFPOSX1_1/a_22_6# 2.40fF
C47 attempt2_4/DFFPOSX1_1/vdd attempt2_4/DFFPOSX1_1/a_22_6# 2.40fF
C48 attempt2_2/DFFPOSX1_0/vdd attempt2_2/DFFPOSX1_0/a_2_6# 4.88fF
C49 attempt2_1/DFFPOSX1_1/vdd attempt2_1/DFFPOSX1_1/a_22_6# 2.40fF
C50 attempt2_3/DFFPOSX1_0/vdd attempt2_3/DFFPOSX1_0/a_34_4# 2.48fF
C51 attempt2_0/DFFPOSX1_0/vdd attempt2_0/DFFPOSX1_0/a_34_4# 2.48fF
C52 attempt2_2/DFFPOSX1_2/vdd attempt2_2/m1_n35_n168# 2.41fF
C53 attempt2_3/DFFPOSX1_2/a_22_6# attempt2_3/DFFPOSX1_2/vdd 2.40fF
C54 attempt2_1/DFFPOSX1_2/vdd attempt2_1/DFFPOSX1_2/a_34_4# 2.48fF
C55 attempt2_3/DFFPOSX1_0/vdd attempt2_3/m1_n29_66# 2.41fF
C56 attempt2_2/DFFPOSX1_0/vdd attempt2_2/DFFPOSX1_0/a_34_4# 2.48fF
C57 attempt2_2/DFFPOSX1_1/vdd attempt2_2/DFFPOSX1_1/a_2_6# 4.88fF
C58 attempt2_1/DFFPOSX1_0/vdd attempt2_1/m1_n29_66# 2.41fF
C59 attempt2_4/m1_n54_n42# attempt2_4/DFFPOSX1_0/vdd 2.20fF
C60 attempt2_3/OR2X1_1/a_2_54# attempt2_3/OR2X1_1/vdd 2.08fF
C61 attempt2_0/DFFPOSX1_1/vdd attempt2_0/DFFPOSX1_1/a_2_6# 4.88fF
C62 attempt2_2/OR2X1_0/vdd attempt2_2/OR2X1_0/a_2_54# 2.08fF
C63 attempt2_4/OR2X1_0/vdd attempt2_4/OR2X1_0/a_2_54# 2.08fF
C64 attempt2_0/OR2X1_0/vdd attempt2_0/OR2X1_0/a_2_54# 2.08fF
C65 attempt2_3/DFFPOSX1_0/vdd attempt2_3/DFFPOSX1_0/a_22_6# 2.40fF
C66 attempt2_0/DFFPOSX1_0/vdd attempt2_0/DFFPOSX1_0/a_22_6# 2.40fF
C67 attempt2_0/DFFPOSX1_1/vdd attempt2_0/DFFPOSX1_1/a_34_4# 2.48fF
C68 attempt2_1/m1_71_n159# attempt2_1/DFFPOSX1_2/vdd 2.20fF
C69 attempt2_4/DFFPOSX1_2/a_22_6# attempt2_4/DFFPOSX1_2/vdd 2.40fF
C70 attempt2_1/DFFPOSX1_2/vdd attempt2_1/DFFPOSX1_2/a_22_6# 2.40fF
C71 attempt2_2/OR2X1_1/vdd attempt2_2/OR2X1_1/a_2_54# 2.08fF
C72 attempt2_0/DFFPOSX1_2/vdd attempt2_0/DFFPOSX1_2/a_2_6# 4.88fF
C73 attempt2_0/m1_n54_n42# attempt2_0/DFFPOSX1_0/vdd 2.20fF
C74 attempt2_3/DFFPOSX1_1/vdd attempt2_3/m1_n31_n51# 2.41fF
C75 attempt2_2/DFFPOSX1_1/vdd attempt2_2/DFFPOSX1_1/a_34_4# 2.48fF
C76 attempt2_1/DFFPOSX1_1/vdd attempt2_1/m1_n31_n51# 2.41fF
C77 attempt2_3/DFFPOSX1_2/vdd attempt2_3/m1_n35_n168# 2.41fF
C78 attempt2_4/DFFPOSX1_2/a_34_4# attempt2_4/DFFPOSX1_2/vdd 2.48fF
C79 attempt2_4/DFFPOSX1_2/vdd attempt2_4/m1_71_n159# 2.20fF
C80 attempt2_3/m1_n54_n42# attempt2_3/DFFPOSX1_0/vdd 2.20fF
C81 attempt2_0/OR2X1_1/vdd attempt2_0/OR2X1_1/a_2_54# 2.08fF
C82 attempt2_3/m1_n64_n214# attempt2_3/DFFPOSX1_1/vdd 2.20fF
C83 attempt2_0/m1_n64_n214# attempt2_0/DFFPOSX1_1/vdd 2.20fF
C84 attempt2_0/DFFPOSX1_1/vdd attempt2_0/DFFPOSX1_1/a_22_6# 2.40fF
C85 attempt2_0/DFFPOSX1_0/gnd Gnd 6.90fF
C86 attempt2_0/DFFPOSX1_0/a_66_6# Gnd 2.10fF
C87 attempt2_0/DFFPOSX1_0/a_2_6# Gnd 2.87fF
C88 attempt2_0/Input1 Gnd 3.01fF
C89 attempt2_0/m1_n29_66# Gnd 5.44fF
C90 attempt2_0/DFFPOSX1_0/vdd Gnd 22.98fF
C91 attempt2_0/DFFPOSX1_1/gnd Gnd 6.90fF
C92 attempt2_0/DFFPOSX1_1/a_66_6# Gnd 2.10fF
C93 attempt2_0/DFFPOSX1_1/a_2_6# Gnd 2.87fF
C94 attempt2_0/m1_n31_n51# Gnd 5.54fF
C95 attempt2_0/DFFPOSX1_1/vdd Gnd 22.98fF
C96 attempt2_0/XOR2X1_0/gnd Gnd 3.69fF
C97 attempt2_0/m1_n64_n214# Gnd 53.33fF
C98 attempt2_0/XOR2X1_0/a_2_6# Gnd 3.28fF
C99 attempt2_0/XOR2X1_0/a_13_43# Gnd 2.84fF
C100 attempt2_0/m1_n54_n42# Gnd 32.43fF
C101 attempt2_0/XOR2X1_0/vdd Gnd 14.77fF
C102 attempt2_0/OR2X1_0/gnd Gnd 2.76fF
C103 attempt2_0/OR2X1_0/a_2_54# Gnd 2.54fF
C104 attempt2_0/m1_133_15# Gnd 3.40fF
C105 attempt2_0/Input3 Gnd 2.30fF
C106 attempt2_0/OR2X1_0/vdd Gnd 9.85fF
C107 attempt2_0/DFFPOSX1_2/gnd Gnd 6.90fF
C108 attempt2_0/DFFPOSX1_2/a_66_6# Gnd 2.10fF
C109 attempt2_0/DFFPOSX1_2/a_2_6# Gnd 2.87fF
C110 attempt2_0/m1_n35_n168# Gnd 5.75fF
C111 attempt2_0/DFFPOSX1_2/vdd Gnd 22.98fF
C112 attempt2_0/XOR2X1_1/gnd Gnd 3.69fF
C113 attempt2_0/m1_71_n159# Gnd 10.24fF
C114 attempt2_0/XOR2X1_1/a_2_6# Gnd 3.28fF
C115 attempt2_0/XOR2X1_1/a_13_43# Gnd 2.84fF
C116 attempt2_0/XOR2X1_1/vdd Gnd 14.77fF
C117 attempt2_0/OR2X1_1/gnd Gnd 2.76fF
C118 attempt2_0/OR2X1_1/a_2_54# Gnd 2.54fF
C119 attempt2_0/OR2X1_1/vdd Gnd 9.85fF
C120 attempt2_1/DFFPOSX1_0/gnd Gnd 6.90fF
C121 attempt2_1/DFFPOSX1_0/a_66_6# Gnd 2.10fF
C122 attempt2_1/DFFPOSX1_0/a_2_6# Gnd 2.87fF
C123 attempt2_1/Input1 Gnd 3.01fF
C124 attempt2_1/m1_n29_66# Gnd 5.44fF
C125 attempt2_1/DFFPOSX1_0/vdd Gnd 22.98fF
C126 attempt2_1/DFFPOSX1_1/gnd Gnd 6.90fF
C127 attempt2_1/DFFPOSX1_1/a_66_6# Gnd 2.10fF
C128 attempt2_1/DFFPOSX1_1/a_2_6# Gnd 2.87fF
C129 attempt2_1/m1_n31_n51# Gnd 5.54fF
C130 attempt2_1/DFFPOSX1_1/vdd Gnd 22.98fF
C131 attempt2_1/XOR2X1_0/gnd Gnd 3.69fF
C132 attempt2_1/m1_n64_n214# Gnd 53.33fF
C133 attempt2_1/XOR2X1_0/a_2_6# Gnd 3.28fF
C134 attempt2_1/XOR2X1_0/a_13_43# Gnd 2.84fF
C135 attempt2_1/m1_n54_n42# Gnd 32.43fF
C136 attempt2_1/XOR2X1_0/vdd Gnd 14.77fF
C137 attempt2_1/OR2X1_0/gnd Gnd 2.76fF
C138 attempt2_1/OR2X1_0/a_2_54# Gnd 2.54fF
C139 attempt2_1/m1_133_15# Gnd 3.40fF
C140 attempt2_1/Input3 Gnd 8.69fF
C141 attempt2_1/OR2X1_0/vdd Gnd 9.85fF
C142 attempt2_1/DFFPOSX1_2/gnd Gnd 6.90fF
C143 attempt2_1/DFFPOSX1_2/a_66_6# Gnd 2.10fF
C144 attempt2_1/DFFPOSX1_2/a_2_6# Gnd 2.87fF
C145 attempt2_1/m1_n35_n168# Gnd 5.75fF
C146 attempt2_1/DFFPOSX1_2/vdd Gnd 22.98fF
C147 attempt2_1/XOR2X1_1/gnd Gnd 3.69fF
C148 attempt2_1/m1_71_n159# Gnd 10.24fF
C149 attempt2_1/XOR2X1_1/a_2_6# Gnd 3.28fF
C150 attempt2_1/XOR2X1_1/a_13_43# Gnd 2.84fF
C151 attempt2_1/XOR2X1_1/vdd Gnd 14.77fF
C152 attempt2_1/OR2X1_1/gnd Gnd 2.76fF
C153 attempt2_1/OR2X1_1/a_2_54# Gnd 2.54fF
C154 attempt2_1/Input2 Gnd 37.23fF
C155 attempt2_1/OR2X1_1/vdd Gnd 9.85fF
C156 attempt2_2/DFFPOSX1_0/gnd Gnd 6.90fF
C157 attempt2_2/DFFPOSX1_0/a_66_6# Gnd 2.10fF
C158 attempt2_2/DFFPOSX1_0/a_2_6# Gnd 2.87fF
C159 attempt2_2/Input1 Gnd 3.01fF
C160 attempt2_2/m1_n29_66# Gnd 5.44fF
C161 attempt2_2/DFFPOSX1_0/vdd Gnd 22.98fF
C162 attempt2_2/DFFPOSX1_1/gnd Gnd 6.90fF
C163 attempt2_2/DFFPOSX1_1/a_66_6# Gnd 2.10fF
C164 attempt2_2/DFFPOSX1_1/a_2_6# Gnd 2.87fF
C165 attempt2_2/m1_n31_n51# Gnd 5.54fF
C166 attempt2_2/DFFPOSX1_1/vdd Gnd 22.98fF
C167 attempt2_2/XOR2X1_0/gnd Gnd 3.69fF
C168 attempt2_2/m1_n64_n214# Gnd 53.33fF
C169 attempt2_2/XOR2X1_0/a_2_6# Gnd 3.28fF
C170 attempt2_2/XOR2X1_0/a_13_43# Gnd 2.84fF
C171 attempt2_2/m1_n54_n42# Gnd 32.43fF
C172 attempt2_2/XOR2X1_0/vdd Gnd 14.77fF
C173 attempt2_2/OR2X1_0/gnd Gnd 2.76fF
C174 attempt2_2/OR2X1_0/a_2_54# Gnd 2.54fF
C175 attempt2_2/m1_133_15# Gnd 3.40fF
C176 attempt2_2/OR2X1_0/vdd Gnd 9.85fF
C177 attempt2_2/DFFPOSX1_2/gnd Gnd 6.90fF
C178 attempt2_2/DFFPOSX1_2/a_66_6# Gnd 2.10fF
C179 attempt2_2/DFFPOSX1_2/a_2_6# Gnd 2.87fF
C180 attempt2_2/m1_n35_n168# Gnd 5.75fF
C181 attempt2_2/DFFPOSX1_2/vdd Gnd 22.98fF
C182 attempt2_2/XOR2X1_1/gnd Gnd 3.69fF
C183 attempt2_2/m1_71_n159# Gnd 10.24fF
C184 attempt2_2/XOR2X1_1/a_2_6# Gnd 3.28fF
C185 attempt2_2/XOR2X1_1/a_13_43# Gnd 2.84fF
C186 attempt2_2/XOR2X1_1/vdd Gnd 14.77fF
C187 attempt2_2/OR2X1_1/gnd Gnd 2.76fF
C188 attempt2_2/OR2X1_1/a_2_54# Gnd 2.54fF
C189 attempt2_2/Input2 Gnd 39.39fF
C190 attempt2_2/OR2X1_1/vdd Gnd 9.85fF
C191 attempt2_3/DFFPOSX1_0/gnd Gnd 6.90fF
C192 attempt2_3/DFFPOSX1_0/a_66_6# Gnd 2.10fF
C193 attempt2_3/DFFPOSX1_0/a_2_6# Gnd 2.87fF
C194 attempt2_3/Input1 Gnd 3.01fF
C195 attempt2_3/m1_n29_66# Gnd 5.44fF
C196 attempt2_3/DFFPOSX1_0/vdd Gnd 22.98fF
C197 attempt2_3/DFFPOSX1_1/gnd Gnd 6.90fF
C198 attempt2_3/DFFPOSX1_1/a_66_6# Gnd 2.10fF
C199 attempt2_3/DFFPOSX1_1/a_2_6# Gnd 2.87fF
C200 attempt2_3/m1_n31_n51# Gnd 5.54fF
C201 attempt2_3/DFFPOSX1_1/vdd Gnd 22.98fF
C202 attempt2_3/XOR2X1_0/gnd Gnd 3.69fF
C203 attempt2_3/m1_n64_n214# Gnd 53.33fF
C204 attempt2_3/XOR2X1_0/a_2_6# Gnd 3.28fF
C205 attempt2_3/XOR2X1_0/a_13_43# Gnd 2.84fF
C206 attempt2_3/m1_n54_n42# Gnd 32.43fF
C207 attempt2_3/XOR2X1_0/vdd Gnd 14.77fF
C208 attempt2_3/OR2X1_0/gnd Gnd 2.76fF
C209 attempt2_3/OR2X1_0/a_2_54# Gnd 2.54fF
C210 attempt2_3/m1_133_15# Gnd 3.40fF
C211 attempt2_3/Input3 Gnd 41.07fF
C212 attempt2_3/OR2X1_0/vdd Gnd 9.85fF
C213 attempt2_3/DFFPOSX1_2/gnd Gnd 6.90fF
C214 attempt2_3/DFFPOSX1_2/a_66_6# Gnd 2.10fF
C215 attempt2_3/DFFPOSX1_2/a_2_6# Gnd 2.87fF
C216 attempt2_3/m1_n35_n168# Gnd 5.75fF
C217 attempt2_3/DFFPOSX1_2/vdd Gnd 22.98fF
C218 attempt2_3/XOR2X1_1/gnd Gnd 3.69fF
C219 attempt2_3/m1_71_n159# Gnd 10.24fF
C220 attempt2_3/XOR2X1_1/a_2_6# Gnd 3.28fF
C221 attempt2_3/XOR2X1_1/a_13_43# Gnd 2.84fF
C222 attempt2_3/XOR2X1_1/vdd Gnd 14.77fF
C223 attempt2_3/OR2X1_1/gnd Gnd 2.76fF
C224 attempt2_3/OR2X1_1/a_2_54# Gnd 2.54fF
C225 attempt2_3/Input2 Gnd 33.76fF
C226 attempt2_3/OR2X1_1/vdd Gnd 9.85fF
C227 attempt2_4/DFFPOSX1_0/gnd Gnd 6.90fF
C228 attempt2_4/DFFPOSX1_0/a_66_6# Gnd 2.10fF
C229 attempt2_4/DFFPOSX1_0/a_2_6# Gnd 2.87fF
C230 attempt2_4/Input1 Gnd 3.01fF
C231 attempt2_4/m1_n29_66# Gnd 5.44fF
C232 attempt2_4/DFFPOSX1_0/vdd Gnd 22.98fF
C233 attempt2_4/DFFPOSX1_1/gnd Gnd 6.90fF
C234 attempt2_4/DFFPOSX1_1/a_66_6# Gnd 2.10fF
C235 attempt2_4/DFFPOSX1_1/a_2_6# Gnd 2.87fF
C236 attempt2_4/m1_n31_n51# Gnd 5.54fF
C237 attempt2_4/DFFPOSX1_1/vdd Gnd 22.98fF
C238 attempt2_4/XOR2X1_0/gnd Gnd 3.69fF
C239 attempt2_4/m1_n64_n214# Gnd 53.33fF
C240 attempt2_4/XOR2X1_0/a_2_6# Gnd 3.28fF
C241 attempt2_4/XOR2X1_0/a_13_43# Gnd 2.84fF
C242 attempt2_4/m1_n54_n42# Gnd 32.43fF
C243 attempt2_4/XOR2X1_0/vdd Gnd 14.77fF
C244 attempt2_4/OR2X1_0/gnd Gnd 2.76fF
C245 attempt2_4/Output1 Gnd 2.78fF
C246 attempt2_4/OR2X1_0/a_2_54# Gnd 2.54fF
C247 attempt2_4/m1_133_15# Gnd 3.40fF
C248 attempt2_4/Input3 Gnd 10.56fF
C249 attempt2_4/OR2X1_0/vdd Gnd 9.85fF
C250 attempt2_4/DFFPOSX1_2/gnd Gnd 6.90fF
C251 attempt2_4/DFFPOSX1_2/a_66_6# Gnd 2.10fF
C252 attempt2_4/DFFPOSX1_2/a_2_6# Gnd 2.87fF
C253 attempt2_4/m1_n35_n168# Gnd 5.75fF
C254 attempt2_4/DFFPOSX1_2/vdd Gnd 22.98fF
C255 attempt2_4/XOR2X1_1/gnd Gnd 3.69fF
C256 attempt2_4/m1_71_n159# Gnd 10.24fF
C257 attempt2_4/XOR2X1_1/a_2_6# Gnd 3.28fF
C258 attempt2_4/XOR2X1_1/a_13_43# Gnd 2.84fF
C259 attempt2_4/XOR2X1_1/vdd Gnd 14.77fF
C260 attempt2_4/OR2X1_1/gnd Gnd 2.76fF
C261 attempt2_4/Output2 Gnd 2.35fF
C262 attempt2_4/OR2X1_1/a_2_54# Gnd 2.54fF
C263 attempt2_4/Input2 Gnd 32.36fF
C264 attempt2_4/OR2X1_1/vdd Gnd 9.85fF
** hspice subcircuit dictionary
.include /home/banturr/Desktop/IntrotoVLSI/Hspice/model_t36s.sp


VDD Vdd Gnd 5V
VIn1 Input1 Gnd PULSE(0 5 0n 0.2n 0.2n 50n 100n)
VIn2 Input2 Gnd PULSE(0 5 0n 0.2n 0.2n 40n 80n)
VIn3 Input3 Gnd PULSE(0 5 0n 0.2n 0.2n 30n 60n)



.options post
.tran 0.01n 60n
.end
